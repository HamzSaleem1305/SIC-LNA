magic
tech sky130A
magscale 1 2
timestamp 1666381508
<< pwell >>
rect -201 -2098 201 2098
<< psubdiff >>
rect -165 2028 -69 2062
rect 69 2028 165 2062
rect -165 1966 -131 2028
rect 131 1966 165 2028
rect -165 -2028 -131 -1966
rect 131 -2028 165 -1966
rect -165 -2062 -69 -2028
rect 69 -2062 165 -2028
<< psubdiffcont >>
rect -69 2028 69 2062
rect -165 -1966 -131 1966
rect 131 -1966 165 1966
rect -69 -2062 69 -2028
<< xpolycontact >>
rect -35 1500 35 1932
rect -35 -1932 35 -1500
<< ppolyres >>
rect -35 -1500 35 1500
<< locali >>
rect -165 2028 -69 2062
rect 69 2028 165 2062
rect -165 1966 -131 2028
rect 131 1966 165 2028
rect -165 -2028 -131 -1966
rect 131 -2028 165 -1966
rect -165 -2062 -69 -2028
rect 69 -2062 165 -2028
<< viali >>
rect -19 1517 19 1914
rect -19 -1914 19 -1517
<< metal1 >>
rect -25 1914 25 1926
rect -25 1517 -19 1914
rect 19 1517 25 1914
rect -25 1505 25 1517
rect -25 -1517 25 -1505
rect -25 -1914 -19 -1517
rect 19 -1914 25 -1517
rect -25 -1926 25 -1914
<< res0p35 >>
rect -37 -1502 37 1502
<< properties >>
string FIXED_BBOX -148 -2045 148 2045
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 15.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 13.815k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
