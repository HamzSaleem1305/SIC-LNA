magic
tech sky130A
magscale 1 2
timestamp 1666418508
<< pwell >>
rect 12980 20580 15600 23390
<< poly >>
rect 14020 23172 14164 23238
rect 15976 21160 16006 21191
rect 14692 21128 14722 21137
rect 14578 21062 14722 21128
rect 15861 21091 16120 21160
<< locali >>
rect 15710 23340 16270 23570
rect 14820 23140 14910 23150
rect 14820 23040 14830 23140
rect 14900 23040 14910 23140
rect 16120 23070 16270 23190
rect 14820 23030 14910 23040
rect 16225 21565 17230 21775
<< viali >>
rect 14830 23040 14900 23140
<< metal1 >>
rect 13650 21780 13800 23385
rect 14090 23180 14740 23240
rect 14041 23132 14111 23151
rect 14041 23050 14050 23132
rect 14102 23050 14111 23132
rect 14041 23031 14111 23050
rect 14241 23132 14311 23151
rect 14241 23050 14250 23132
rect 14302 23050 14311 23132
rect 14241 23031 14311 23050
rect 14431 23132 14501 23151
rect 14431 23050 14440 23132
rect 14492 23050 14501 23132
rect 14431 23031 14501 23050
rect 14621 23132 14691 23151
rect 14621 23050 14630 23132
rect 14682 23050 14691 23132
rect 14621 23031 14691 23050
rect 14810 23140 14920 23160
rect 14810 23040 14830 23140
rect 14900 23040 14920 23140
rect 14810 23020 14920 23040
rect 15260 22760 15420 23480
rect 15950 23230 16030 23280
rect 15901 23172 15971 23191
rect 15901 23090 15910 23172
rect 15962 23090 15971 23172
rect 15901 23071 15971 23090
rect 16091 23172 16161 23191
rect 16091 23090 16100 23172
rect 16152 23090 16161 23172
rect 16091 23071 16161 23090
rect 13480 21630 13800 21780
rect 13000 21070 13560 21190
rect 13710 21120 13800 21630
rect 15801 21292 15871 21311
rect 13951 21252 14021 21271
rect 13951 21170 13960 21252
rect 14012 21170 14021 21252
rect 13951 21151 14021 21170
rect 14141 21252 14211 21271
rect 14141 21170 14150 21252
rect 14202 21170 14211 21252
rect 14141 21151 14211 21170
rect 14331 21252 14401 21271
rect 14331 21170 14340 21252
rect 14392 21170 14401 21252
rect 14331 21151 14401 21170
rect 14521 21252 14591 21271
rect 14521 21170 14530 21252
rect 14582 21170 14591 21252
rect 14521 21151 14591 21170
rect 14721 21252 14791 21271
rect 14721 21170 14730 21252
rect 14782 21170 14791 21252
rect 14721 21151 14791 21170
rect 15290 21150 15390 21290
rect 15801 21210 15810 21292
rect 15862 21210 15871 21292
rect 15801 21191 15871 21210
rect 16001 21292 16071 21311
rect 16001 21210 16010 21292
rect 16062 21210 16071 21292
rect 16001 21191 16071 21210
rect 13000 16224 13120 21070
rect 13710 21040 14650 21120
rect 15290 21080 16120 21150
rect 13000 16104 13810 16224
<< via1 >>
rect 14050 23050 14102 23132
rect 14250 23050 14302 23132
rect 14440 23050 14492 23132
rect 14630 23050 14682 23132
rect 14830 23040 14900 23140
rect 15910 23090 15962 23172
rect 16100 23090 16152 23172
rect 13960 21170 14012 21252
rect 14150 21170 14202 21252
rect 14340 21170 14392 21252
rect 14530 21170 14582 21252
rect 14730 21170 14782 21252
rect 15810 21210 15862 21292
rect 16010 21210 16062 21292
<< metal2 >>
rect 15901 23190 15971 23191
rect 16091 23190 16161 23191
rect 15901 23172 16161 23190
rect 14041 23150 14111 23151
rect 14241 23150 14311 23151
rect 14431 23150 14501 23151
rect 14621 23150 14691 23151
rect 14041 23140 14910 23150
rect 14041 23132 14830 23140
rect 14041 23050 14050 23132
rect 14102 23050 14250 23132
rect 14302 23050 14440 23132
rect 14492 23050 14630 23132
rect 14682 23050 14830 23132
rect 14041 23040 14830 23050
rect 14900 23040 14910 23140
rect 15901 23090 15910 23172
rect 15962 23090 16100 23172
rect 16152 23090 16161 23172
rect 15901 23071 16161 23090
rect 15920 23070 16160 23071
rect 14041 23031 14910 23040
rect 14060 23030 14910 23031
rect 15801 21310 15871 21311
rect 16001 21310 16071 21311
rect 15801 21292 16071 21310
rect 15801 21274 15810 21292
rect 13964 21271 15810 21274
rect 13951 21252 15810 21271
rect 13951 21170 13960 21252
rect 14012 21170 14150 21252
rect 14202 21170 14340 21252
rect 14392 21170 14530 21252
rect 14582 21170 14730 21252
rect 14782 21210 15810 21252
rect 15862 21210 16010 21292
rect 16062 21274 16071 21292
rect 16062 21210 16074 21274
rect 14782 21170 16074 21210
rect 13951 21151 16074 21170
rect 13964 21146 16074 21151
rect 15615 20310 15745 21146
use sky130_fd_pr__pfet_01v8_XGJ6MR  XM19
timestamp 1666417074
transform 1 0 15991 0 1 22189
box -311 -1219 311 1219
use sky130_fd_pr__nfet_01v8_lvt_CULS5R  XM22
timestamp 1666417074
transform 1 0 14371 0 1 22150
box -551 -1210 551 1210
use sky130_fd_pr__res_high_po_0p35_S8HYGH  XR13
timestamp 1666417074
transform 1 0 15341 0 1 22178
box -201 -1218 201 1218
use sky130_fd_pr__res_high_po_0p35_SVGS7M  XR18
timestamp 1666417074
transform 1 0 13521 0 1 21588
box -201 -648 201 648
use partition3  partition3_0
timestamp 1666417074
transform 1 0 9850 0 1 21340
box -3860 -11100 15212 3114
<< labels >>
flabel metal1 15330 23430 15330 23430 0 FreeSans 1600 0 0 0 VB0_6
flabel metal1 13710 23310 13710 23310 0 FreeSans 1600 0 0 0 VSI2
flabel locali 16150 23460 16150 23460 0 FreeSans 1600 0 0 0 VDD
flabel metal2 15010 21210 15010 21210 0 FreeSans 1600 0 0 0 Vo2
flabel via1 14870 23090 14870 23090 0 FreeSans 1600 0 0 0 VSS
<< end >>
