magic
tech sky130A
timestamp 1640952342
<< error_p >>
rect -54 -250 -25 250
rect 25 -250 54 250
<< nmos >>
rect -25 -250 25 250
<< ndiff >>
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
<< ndiffc >>
rect -48 -244 -31 244
rect 31 -244 48 244
<< poly >>
rect -25 250 25 263
rect -25 -263 25 -250
<< locali >>
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
<< viali >>
rect -48 -244 -31 244
rect 31 -244 48 244
<< metal1 >>
rect -51 244 -28 250
rect -51 -244 -48 244
rect -31 -244 -28 244
rect -51 -250 -28 -244
rect 28 244 51 250
rect 28 -244 31 244
rect 48 -244 51 244
rect 28 -250 51 -244
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
