magic
tech sky130A
magscale 1 2
timestamp 1666381508
<< error_p >>
rect -221 715 -163 721
rect -29 715 29 721
rect 163 715 221 721
rect -221 681 -209 715
rect -29 681 -17 715
rect 163 681 175 715
rect -221 675 -163 681
rect -29 675 29 681
rect 163 675 221 681
rect -317 -681 -259 -675
rect -125 -681 -67 -675
rect 67 -681 125 -675
rect 259 -681 317 -675
rect -317 -715 -305 -681
rect -125 -715 -113 -681
rect 67 -715 79 -681
rect 259 -715 271 -681
rect -317 -721 -259 -715
rect -125 -721 -67 -715
rect 67 -721 125 -715
rect 259 -721 317 -715
<< pwell >>
rect -503 -853 503 853
<< nmoslvt >>
rect -303 -643 -273 643
rect -207 -643 -177 643
rect -111 -643 -81 643
rect -15 -643 15 643
rect 81 -643 111 643
rect 177 -643 207 643
rect 273 -643 303 643
<< ndiff >>
rect -365 631 -303 643
rect -365 -631 -353 631
rect -319 -631 -303 631
rect -365 -643 -303 -631
rect -273 631 -207 643
rect -273 -631 -257 631
rect -223 -631 -207 631
rect -273 -643 -207 -631
rect -177 631 -111 643
rect -177 -631 -161 631
rect -127 -631 -111 631
rect -177 -643 -111 -631
rect -81 631 -15 643
rect -81 -631 -65 631
rect -31 -631 -15 631
rect -81 -643 -15 -631
rect 15 631 81 643
rect 15 -631 31 631
rect 65 -631 81 631
rect 15 -643 81 -631
rect 111 631 177 643
rect 111 -631 127 631
rect 161 -631 177 631
rect 111 -643 177 -631
rect 207 631 273 643
rect 207 -631 223 631
rect 257 -631 273 631
rect 207 -643 273 -631
rect 303 631 365 643
rect 303 -631 319 631
rect 353 -631 365 631
rect 303 -643 365 -631
<< ndiffc >>
rect -353 -631 -319 631
rect -257 -631 -223 631
rect -161 -631 -127 631
rect -65 -631 -31 631
rect 31 -631 65 631
rect 127 -631 161 631
rect 223 -631 257 631
rect 319 -631 353 631
<< psubdiff >>
rect -467 783 -371 817
rect 371 783 467 817
rect -467 721 -433 783
rect 433 721 467 783
rect -467 -783 -433 -721
rect 433 -783 467 -721
rect -467 -817 -371 -783
rect 371 -817 467 -783
<< psubdiffcont >>
rect -371 783 371 817
rect -467 -721 -433 721
rect 433 -721 467 721
rect -371 -817 371 -783
<< poly >>
rect -225 715 -159 731
rect -225 681 -209 715
rect -175 681 -159 715
rect -303 643 -273 669
rect -225 665 -159 681
rect -33 715 33 731
rect -33 681 -17 715
rect 17 681 33 715
rect -207 643 -177 665
rect -111 643 -81 669
rect -33 665 33 681
rect 159 715 225 731
rect 159 681 175 715
rect 209 681 225 715
rect -15 643 15 665
rect 81 643 111 669
rect 159 665 225 681
rect 177 643 207 665
rect 273 643 303 669
rect -303 -665 -273 -643
rect -321 -681 -255 -665
rect -207 -669 -177 -643
rect -111 -665 -81 -643
rect -321 -715 -305 -681
rect -271 -715 -255 -681
rect -321 -731 -255 -715
rect -129 -681 -63 -665
rect -15 -669 15 -643
rect 81 -665 111 -643
rect -129 -715 -113 -681
rect -79 -715 -63 -681
rect -129 -731 -63 -715
rect 63 -681 129 -665
rect 177 -669 207 -643
rect 273 -665 303 -643
rect 63 -715 79 -681
rect 113 -715 129 -681
rect 63 -731 129 -715
rect 255 -681 321 -665
rect 255 -715 271 -681
rect 305 -715 321 -681
rect 255 -731 321 -715
<< polycont >>
rect -209 681 -175 715
rect -17 681 17 715
rect 175 681 209 715
rect -305 -715 -271 -681
rect -113 -715 -79 -681
rect 79 -715 113 -681
rect 271 -715 305 -681
<< locali >>
rect -467 783 -371 817
rect 371 783 467 817
rect -467 721 -433 783
rect 433 721 467 783
rect -225 681 -209 715
rect -175 681 -159 715
rect -33 681 -17 715
rect 17 681 33 715
rect 159 681 175 715
rect 209 681 225 715
rect -353 631 -319 647
rect -353 -647 -319 -631
rect -257 631 -223 647
rect -257 -647 -223 -631
rect -161 631 -127 647
rect -161 -647 -127 -631
rect -65 631 -31 647
rect -65 -647 -31 -631
rect 31 631 65 647
rect 31 -647 65 -631
rect 127 631 161 647
rect 127 -647 161 -631
rect 223 631 257 647
rect 223 -647 257 -631
rect 319 631 353 647
rect 319 -647 353 -631
rect -321 -715 -305 -681
rect -271 -715 -255 -681
rect -129 -715 -113 -681
rect -79 -715 -63 -681
rect 63 -715 79 -681
rect 113 -715 129 -681
rect 255 -715 271 -681
rect 305 -715 321 -681
rect -467 -783 -433 -721
rect 433 -783 467 -721
rect -467 -817 -371 -783
rect 371 -817 467 -783
<< viali >>
rect -209 681 -175 715
rect -17 681 17 715
rect 175 681 209 715
rect -353 -631 -319 631
rect -257 -631 -223 631
rect -161 -631 -127 631
rect -65 -631 -31 631
rect 31 -631 65 631
rect 127 -631 161 631
rect 223 -631 257 631
rect 319 -631 353 631
rect -305 -715 -271 -681
rect -113 -715 -79 -681
rect 79 -715 113 -681
rect 271 -715 305 -681
<< metal1 >>
rect -221 715 -163 721
rect -221 681 -209 715
rect -175 681 -163 715
rect -221 675 -163 681
rect -29 715 29 721
rect -29 681 -17 715
rect 17 681 29 715
rect -29 675 29 681
rect 163 715 221 721
rect 163 681 175 715
rect 209 681 221 715
rect 163 675 221 681
rect -359 631 -313 643
rect -359 -631 -353 631
rect -319 -631 -313 631
rect -359 -643 -313 -631
rect -263 631 -217 643
rect -263 -631 -257 631
rect -223 -631 -217 631
rect -263 -643 -217 -631
rect -167 631 -121 643
rect -167 -631 -161 631
rect -127 -631 -121 631
rect -167 -643 -121 -631
rect -71 631 -25 643
rect -71 -631 -65 631
rect -31 -631 -25 631
rect -71 -643 -25 -631
rect 25 631 71 643
rect 25 -631 31 631
rect 65 -631 71 631
rect 25 -643 71 -631
rect 121 631 167 643
rect 121 -631 127 631
rect 161 -631 167 631
rect 121 -643 167 -631
rect 217 631 263 643
rect 217 -631 223 631
rect 257 -631 263 631
rect 217 -643 263 -631
rect 313 631 359 643
rect 313 -631 319 631
rect 353 -631 359 631
rect 313 -643 359 -631
rect -317 -681 -259 -675
rect -317 -715 -305 -681
rect -271 -715 -259 -681
rect -317 -721 -259 -715
rect -125 -681 -67 -675
rect -125 -715 -113 -681
rect -79 -715 -67 -681
rect -125 -721 -67 -715
rect 67 -681 125 -675
rect 67 -715 79 -681
rect 113 -715 125 -681
rect 67 -721 125 -715
rect 259 -681 317 -675
rect 259 -715 271 -681
rect 305 -715 317 -681
rect 259 -721 317 -715
<< properties >>
string FIXED_BBOX -450 -800 450 800
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 6.428571428571429 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
