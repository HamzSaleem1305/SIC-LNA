magic
tech sky130A
magscale 1 2
timestamp 1666367785
<< error_p >>
rect -269 1072 -211 1078
rect -77 1072 -19 1078
rect 115 1072 173 1078
rect 307 1072 365 1078
rect -269 1038 -257 1072
rect -77 1038 -65 1072
rect 115 1038 127 1072
rect 307 1038 319 1072
rect -269 1032 -211 1038
rect -77 1032 -19 1038
rect 115 1032 173 1038
rect 307 1032 365 1038
rect -365 -1038 -307 -1032
rect -173 -1038 -115 -1032
rect 19 -1038 77 -1032
rect 211 -1038 269 -1032
rect -365 -1072 -353 -1038
rect -173 -1072 -161 -1038
rect 19 -1072 31 -1038
rect 211 -1072 223 -1038
rect -365 -1078 -307 -1072
rect -173 -1078 -115 -1072
rect 19 -1078 77 -1072
rect 211 -1078 269 -1072
<< pwell >>
rect -551 -1210 551 1210
<< nmoslvt >>
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
<< ndiff >>
rect -413 988 -351 1000
rect -413 -988 -401 988
rect -367 -988 -351 988
rect -413 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 413 1000
rect 351 -988 367 988
rect 401 -988 413 988
rect 351 -1000 413 -988
<< ndiffc >>
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
<< psubdiff >>
rect -515 1140 -419 1174
rect 419 1140 515 1174
rect -515 1078 -481 1140
rect 481 1078 515 1140
rect -515 -1140 -481 -1078
rect 481 -1140 515 -1078
rect -515 -1174 -419 -1140
rect 419 -1174 515 -1140
<< psubdiffcont >>
rect -419 1140 419 1174
rect -515 -1078 -481 1078
rect 481 -1078 515 1078
rect -419 -1174 419 -1140
<< poly >>
rect -273 1072 -207 1088
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -351 1000 -321 1026
rect -273 1022 -207 1038
rect -81 1072 -15 1088
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect -255 1000 -225 1022
rect -159 1000 -129 1026
rect -81 1022 -15 1038
rect 111 1072 177 1088
rect 111 1038 127 1072
rect 161 1038 177 1072
rect -63 1000 -33 1022
rect 33 1000 63 1026
rect 111 1022 177 1038
rect 303 1072 369 1088
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 129 1000 159 1022
rect 225 1000 255 1026
rect 303 1022 369 1038
rect 321 1000 351 1022
rect -351 -1022 -321 -1000
rect -369 -1038 -303 -1022
rect -255 -1026 -225 -1000
rect -159 -1022 -129 -1000
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -369 -1088 -303 -1072
rect -177 -1038 -111 -1022
rect -63 -1026 -33 -1000
rect 33 -1022 63 -1000
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect -177 -1088 -111 -1072
rect 15 -1038 81 -1022
rect 129 -1026 159 -1000
rect 225 -1022 255 -1000
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 15 -1088 81 -1072
rect 207 -1038 273 -1022
rect 321 -1026 351 -1000
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 207 -1088 273 -1072
<< polycont >>
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
<< locali >>
rect -515 1140 -419 1174
rect 419 1140 515 1174
rect -515 1078 -481 1140
rect 481 1078 515 1140
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect 111 1038 127 1072
rect 161 1038 177 1072
rect 303 1038 319 1072
rect 353 1038 369 1072
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect -515 -1140 -481 -1078
rect 481 -1140 515 -1078
rect -515 -1174 -419 -1140
rect 419 -1174 515 -1140
<< viali >>
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
<< metal1 >>
rect -269 1072 -211 1078
rect -269 1038 -257 1072
rect -223 1038 -211 1072
rect -269 1032 -211 1038
rect -77 1072 -19 1078
rect -77 1038 -65 1072
rect -31 1038 -19 1072
rect -77 1032 -19 1038
rect 115 1072 173 1078
rect 115 1038 127 1072
rect 161 1038 173 1072
rect 115 1032 173 1038
rect 307 1072 365 1078
rect 307 1038 319 1072
rect 353 1038 365 1072
rect 307 1032 365 1038
rect -407 988 -361 1000
rect -407 -988 -401 988
rect -367 -988 -361 988
rect -407 -1000 -361 -988
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect 361 988 407 1000
rect 361 -988 367 988
rect 401 -988 407 988
rect 361 -1000 407 -988
rect -365 -1038 -307 -1032
rect -365 -1072 -353 -1038
rect -319 -1072 -307 -1038
rect -365 -1078 -307 -1072
rect -173 -1038 -115 -1032
rect -173 -1072 -161 -1038
rect -127 -1072 -115 -1038
rect -173 -1078 -115 -1072
rect 19 -1038 77 -1032
rect 19 -1072 31 -1038
rect 65 -1072 77 -1038
rect 19 -1078 77 -1072
rect 211 -1038 269 -1032
rect 211 -1072 223 -1038
rect 257 -1072 269 -1038
rect 211 -1078 269 -1072
<< properties >>
string FIXED_BBOX -498 -1157 498 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
