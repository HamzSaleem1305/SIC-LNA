magic
tech sky130A
magscale 1 2
timestamp 1666373124
<< pwell >>
rect 1282 210 6247 3375
<< psubdiff >>
rect 1372 3247 6168 3266
rect 1372 3164 1611 3247
rect 5894 3164 6168 3247
rect 1372 3131 6168 3164
rect 1372 3100 1507 3131
rect 1372 466 1401 3100
rect 1474 466 1507 3100
rect 6026 3109 6168 3131
rect 1372 414 1507 466
rect 6026 475 6064 3109
rect 6137 475 6168 3109
rect 6026 414 6168 475
rect 1372 394 6168 414
rect 1372 311 1653 394
rect 5936 311 6168 394
rect 1372 286 6168 311
<< psubdiffcont >>
rect 1611 3164 5894 3247
rect 1401 466 1474 3100
rect 6064 475 6137 3109
rect 1653 311 5936 394
<< poly >>
rect 2770 5600 2920 5670
rect 5440 5645 5662 5716
rect 2770 5590 2800 5600
rect 1896 5172 1964 5230
rect 3442 3558 3472 3569
rect 3328 3492 3472 3558
rect 5422 3522 5680 3593
rect 5298 2989 5416 3010
rect 5298 2949 5319 2989
rect 5391 2949 5416 2989
rect 5298 2930 5416 2949
rect 1778 2871 1869 2891
rect 1778 2809 1798 2871
rect 1850 2851 1869 2871
rect 1973 2853 2048 2871
rect 1850 2809 1896 2851
rect 1973 2848 1987 2853
rect 1778 2772 1896 2809
rect 1954 2807 1987 2848
rect 2034 2848 2048 2853
rect 2327 2849 2402 2867
rect 2034 2807 2072 2848
rect 2327 2846 2341 2849
rect 1954 2791 2072 2807
rect 1954 2746 1984 2791
rect 2042 2748 2072 2791
rect 2306 2803 2341 2846
rect 2388 2846 2402 2849
rect 2680 2848 2755 2865
rect 3033 2848 3108 2866
rect 3384 2848 3459 2866
rect 3738 2849 3813 2867
rect 4088 2849 4163 2866
rect 3738 2848 3752 2849
rect 2658 2847 2776 2848
rect 2388 2803 2424 2846
rect 2306 2787 2424 2803
rect 2306 2744 2336 2787
rect 2394 2746 2424 2787
rect 2658 2801 2694 2847
rect 2741 2801 2776 2847
rect 2658 2785 2776 2801
rect 2658 2746 2688 2785
rect 2746 2748 2776 2785
rect 3010 2802 3047 2848
rect 3094 2802 3128 2848
rect 3010 2786 3128 2802
rect 3010 2746 3040 2786
rect 3098 2748 3128 2786
rect 3362 2802 3398 2848
rect 3445 2802 3480 2848
rect 3362 2786 3480 2802
rect 3362 2746 3392 2786
rect 3450 2748 3480 2786
rect 3714 2803 3752 2848
rect 3799 2848 3813 2849
rect 4066 2848 4184 2849
rect 4440 2848 4515 2865
rect 4793 2848 4868 2865
rect 5142 2848 5217 2865
rect 3799 2803 3832 2848
rect 3714 2787 3832 2803
rect 3714 2746 3744 2787
rect 3802 2748 3832 2787
rect 4066 2802 4102 2848
rect 4149 2802 4184 2848
rect 4066 2786 4184 2802
rect 4066 2747 4096 2786
rect 4154 2749 4184 2786
rect 4418 2847 4536 2848
rect 4418 2801 4454 2847
rect 4501 2801 4536 2847
rect 4418 2785 4536 2801
rect 4418 2746 4448 2785
rect 4506 2748 4536 2785
rect 4770 2847 4888 2848
rect 4770 2801 4807 2847
rect 4854 2801 4888 2847
rect 4770 2785 4888 2801
rect 4770 2746 4800 2785
rect 4858 2748 4888 2785
rect 5122 2847 5240 2848
rect 5122 2801 5156 2847
rect 5203 2801 5240 2847
rect 5122 2785 5240 2801
rect 5122 2746 5152 2785
rect 5210 2748 5240 2785
rect 5298 2772 5328 2930
rect 5386 2772 5416 2930
rect 5496 2849 5571 2865
rect 5474 2847 5592 2849
rect 5474 2801 5510 2847
rect 5557 2801 5592 2847
rect 5669 2847 5744 2865
rect 5669 2840 5683 2847
rect 5474 2785 5592 2801
rect 5474 2747 5504 2785
rect 5562 2749 5592 2785
rect 5650 2801 5683 2840
rect 5730 2840 5744 2847
rect 5730 2801 5768 2840
rect 5650 2785 5768 2801
rect 5650 2762 5680 2785
rect 5738 2744 5768 2785
rect 1778 696 1808 748
rect 1866 696 1896 744
rect 1778 678 1896 696
rect 1778 646 1809 678
rect 1795 632 1809 646
rect 1856 646 1896 678
rect 2130 690 2160 747
rect 2218 690 2248 745
rect 2130 672 2248 690
rect 1856 632 1870 646
rect 2130 645 2159 672
rect 1795 616 1870 632
rect 2145 626 2159 645
rect 2206 645 2248 672
rect 2482 693 2512 747
rect 2570 693 2600 745
rect 2482 675 2600 693
rect 2482 645 2517 675
rect 2206 626 2220 645
rect 2145 610 2220 626
rect 2503 629 2517 645
rect 2564 645 2600 675
rect 2834 693 2864 747
rect 2922 693 2952 745
rect 2834 675 2952 693
rect 2834 645 2865 675
rect 2564 629 2578 645
rect 2503 613 2578 629
rect 2851 629 2865 645
rect 2912 645 2952 675
rect 3186 693 3216 748
rect 3274 693 3304 746
rect 3186 675 3304 693
rect 3186 646 3216 675
rect 2912 629 2926 645
rect 2851 613 2926 629
rect 3202 629 3216 646
rect 3263 646 3304 675
rect 3538 692 3568 748
rect 3626 692 3656 746
rect 3538 674 3656 692
rect 3538 646 3567 674
rect 3263 629 3277 646
rect 3202 613 3277 629
rect 3553 628 3567 646
rect 3614 646 3656 674
rect 3890 690 3920 749
rect 3978 690 4008 747
rect 3890 672 4008 690
rect 3890 647 3918 672
rect 3614 628 3628 646
rect 3553 612 3628 628
rect 3904 626 3918 647
rect 3965 647 4008 672
rect 4242 693 4272 749
rect 4330 693 4360 747
rect 4242 675 4360 693
rect 4242 647 4273 675
rect 3965 626 3979 647
rect 3904 610 3979 626
rect 4259 629 4273 647
rect 4320 647 4360 675
rect 4594 689 4624 749
rect 4682 689 4712 747
rect 4594 671 4712 689
rect 4594 647 4623 671
rect 4320 629 4334 647
rect 4259 613 4334 629
rect 4609 625 4623 647
rect 4670 647 4712 671
rect 4946 691 4976 748
rect 5034 691 5064 746
rect 4946 673 5064 691
rect 4670 625 4684 647
rect 4946 646 4977 673
rect 4609 609 4684 625
rect 4963 627 4977 646
rect 5024 646 5064 673
rect 5298 689 5328 749
rect 5386 689 5416 747
rect 5298 671 5416 689
rect 5298 647 5327 671
rect 5024 627 5038 646
rect 4963 611 5038 627
rect 5313 625 5327 647
rect 5374 647 5416 671
rect 5650 700 5680 750
rect 5738 700 5768 748
rect 5650 670 5770 700
rect 5374 625 5388 647
rect 5313 609 5388 625
rect 5650 590 5670 670
rect 5750 590 5770 670
rect 5650 560 5770 590
<< polycont >>
rect 5319 2949 5391 2989
rect 1798 2809 1850 2871
rect 1987 2807 2034 2853
rect 2341 2803 2388 2849
rect 2694 2801 2741 2847
rect 3047 2802 3094 2848
rect 3398 2802 3445 2848
rect 3752 2803 3799 2849
rect 4102 2802 4149 2848
rect 4454 2801 4501 2847
rect 4807 2801 4854 2847
rect 5156 2801 5203 2847
rect 5510 2801 5557 2847
rect 5683 2801 5730 2847
rect 1809 632 1856 678
rect 2159 626 2206 672
rect 2517 629 2564 675
rect 2865 629 2912 675
rect 3216 629 3263 675
rect 3567 628 3614 674
rect 3918 626 3965 672
rect 4273 629 4320 675
rect 4623 625 4670 671
rect 4977 627 5024 673
rect 5327 625 5374 671
rect 5670 590 5750 670
<< locali >>
rect 5239 5769 5859 5921
rect 5676 5500 5828 5619
rect 1957 5003 2106 5139
rect 1372 3247 6168 3266
rect 1372 3164 1611 3247
rect 5894 3164 6168 3247
rect 1372 3131 6168 3164
rect 1372 3100 1507 3131
rect 1372 466 1401 3100
rect 1474 466 1507 3100
rect 6026 3109 6168 3131
rect 4420 3020 4540 3030
rect 4420 2960 4430 3020
rect 4530 2960 4540 3020
rect 1778 2871 1869 2891
rect 4420 2874 4540 2960
rect 5298 2989 5416 3010
rect 5298 2949 5319 2989
rect 5391 2949 5416 2989
rect 5298 2930 5416 2949
rect 1778 2809 1798 2871
rect 1850 2809 1869 2871
rect 1778 2791 1869 2809
rect 1912 2853 5772 2874
rect 1912 2807 1987 2853
rect 2034 2849 5772 2853
rect 2034 2807 2341 2849
rect 1912 2803 2341 2807
rect 2388 2848 3752 2849
rect 2388 2847 3047 2848
rect 2388 2803 2694 2847
rect 1912 2801 2694 2803
rect 2741 2802 3047 2847
rect 3094 2802 3398 2848
rect 3445 2803 3752 2848
rect 3799 2848 5772 2849
rect 3799 2803 4102 2848
rect 3445 2802 4102 2803
rect 4149 2847 5772 2848
rect 4149 2802 4454 2847
rect 2741 2801 4454 2802
rect 4501 2801 4807 2847
rect 4854 2801 5156 2847
rect 5203 2801 5510 2847
rect 5557 2801 5683 2847
rect 5730 2801 5772 2847
rect 1912 2795 5772 2801
rect 1973 2791 2048 2795
rect 2327 2787 2402 2795
rect 2680 2785 2755 2795
rect 3033 2786 3108 2795
rect 3384 2786 3459 2795
rect 3738 2787 3813 2795
rect 4088 2786 4163 2795
rect 4420 2790 4540 2795
rect 4440 2785 4515 2790
rect 4793 2785 4868 2795
rect 5142 2785 5217 2795
rect 5496 2785 5571 2795
rect 5669 2785 5744 2795
rect 1795 678 1870 696
rect 1795 676 1809 678
rect 1765 632 1809 676
rect 1856 676 1870 678
rect 2145 676 2220 690
rect 2503 676 2578 693
rect 2851 676 2926 693
rect 3202 676 3277 693
rect 3553 676 3628 692
rect 3904 676 3979 690
rect 4259 676 4334 693
rect 4609 676 4684 689
rect 4963 676 5038 691
rect 5313 676 5388 689
rect 1856 675 5456 676
rect 1856 672 2517 675
rect 1856 632 2159 672
rect 1765 626 2159 632
rect 2206 629 2517 672
rect 2564 629 2865 675
rect 2912 629 3216 675
rect 3263 674 4273 675
rect 3263 629 3567 674
rect 2206 628 3567 629
rect 3614 672 4273 674
rect 3614 628 3918 672
rect 2206 626 3918 628
rect 3965 629 4273 672
rect 4320 673 5456 675
rect 4320 671 4977 673
rect 4320 629 4623 671
rect 3965 626 4623 629
rect 1765 625 4623 626
rect 4670 627 4977 671
rect 5024 671 5456 673
rect 5024 627 5327 671
rect 4670 625 5327 627
rect 5374 625 5456 671
rect 1765 607 5456 625
rect 5650 670 5770 700
rect 1765 550 1895 607
rect 5650 590 5670 670
rect 5750 590 5770 670
rect 5650 570 5770 590
rect 1765 491 1780 550
rect 1879 491 1895 550
rect 1765 480 1895 491
rect 5640 550 5780 570
rect 1372 414 1507 466
rect 5640 460 5660 550
rect 5760 460 5780 550
rect 5640 450 5780 460
rect 6026 475 6064 3109
rect 6137 475 6168 3109
rect 6026 414 6168 475
rect 1372 394 6168 414
rect 1372 311 1653 394
rect 5936 311 6168 394
rect 1372 286 6168 311
rect 2159 -84 5303 286
<< viali >>
rect 4430 2960 4530 3020
rect 5319 2949 5391 2989
rect 1798 2809 1850 2871
rect 1780 491 1879 550
rect 5660 460 5760 550
rect 2800 330 2980 390
<< metal1 >>
rect 1870 5780 4540 5900
rect 1870 5170 1990 5780
rect 3040 5680 3140 5690
rect 3040 5660 3050 5680
rect 2850 5620 3050 5660
rect 3130 5660 3140 5680
rect 3130 5620 3490 5660
rect 2850 5610 3490 5620
rect 2791 5570 2861 5580
rect 2791 5470 2800 5570
rect 2852 5470 2861 5570
rect 2791 5460 2861 5470
rect 2991 5570 3061 5580
rect 2991 5470 3000 5570
rect 3052 5470 3061 5570
rect 2991 5460 3061 5470
rect 3181 5570 3251 5580
rect 3181 5470 3190 5570
rect 3242 5470 3251 5570
rect 3181 5460 3251 5470
rect 3371 5570 3441 5580
rect 3371 5470 3380 5570
rect 3432 5470 3441 5570
rect 3371 5460 3441 5470
rect 4420 5200 4540 5780
rect 5510 5660 5590 5720
rect 5471 5610 5541 5620
rect 5471 5510 5480 5610
rect 5532 5510 5541 5610
rect 5471 5500 5541 5510
rect 5661 5610 5731 5620
rect 5661 5510 5670 5610
rect 5722 5510 5731 5610
rect 5661 5500 5731 5510
rect 2711 3700 2781 3710
rect 1778 2871 1870 3696
rect 2711 3600 2720 3700
rect 2772 3600 2781 3700
rect 2711 3590 2781 3600
rect 2891 3700 2961 3710
rect 2891 3600 2900 3700
rect 2952 3600 2961 3700
rect 2891 3590 2961 3600
rect 3081 3700 3151 3710
rect 3081 3600 3090 3700
rect 3142 3600 3151 3700
rect 3081 3590 3151 3600
rect 3271 3700 3341 3710
rect 3271 3600 3280 3700
rect 3332 3600 3341 3700
rect 3271 3590 3341 3600
rect 3461 3700 3531 3710
rect 3461 3600 3470 3700
rect 3522 3600 3531 3700
rect 3461 3590 3531 3600
rect 1898 3540 1966 3547
rect 1898 3489 1909 3540
rect 1899 3479 1909 3489
rect 1961 3479 1966 3540
rect 2750 3500 3390 3550
rect 1899 3470 1966 3479
rect 4420 3030 4540 3990
rect 5371 3730 5441 3740
rect 5371 3630 5380 3730
rect 5432 3630 5441 3730
rect 5371 3620 5441 3630
rect 5571 3730 5641 3740
rect 5571 3630 5580 3730
rect 5632 3630 5641 3730
rect 5571 3620 5641 3630
rect 5420 3589 5680 3590
rect 5298 3471 5683 3589
rect 4410 3020 4550 3030
rect 4410 2960 4430 3020
rect 4530 2960 4550 3020
rect 4410 2940 4550 2960
rect 5298 2989 5416 3471
rect 5298 2949 5319 2989
rect 5391 2949 5416 2989
rect 5298 2930 5416 2949
rect 1778 2809 1798 2871
rect 1850 2809 1870 2871
rect 1778 2792 1870 2809
rect 1901 2849 2122 2895
rect 1778 2791 1869 2792
rect 1806 2728 1868 2738
rect 1806 2636 1810 2728
rect 1864 2636 1868 2728
rect 1901 2727 1947 2849
rect 1976 2731 2041 2744
rect 1806 2626 1868 2636
rect 1976 2642 1983 2731
rect 2035 2642 2041 2731
rect 2076 2718 2122 2849
rect 2257 2846 2478 2892
rect 2154 2728 2216 2738
rect 1976 2630 2041 2642
rect 2154 2636 2158 2728
rect 2212 2636 2216 2728
rect 2257 2724 2303 2846
rect 2333 2733 2398 2746
rect 2154 2626 2216 2636
rect 2333 2644 2340 2733
rect 2392 2644 2398 2733
rect 2432 2715 2478 2846
rect 2610 2851 2831 2897
rect 2510 2734 2572 2744
rect 2333 2632 2398 2644
rect 2510 2642 2514 2734
rect 2568 2642 2572 2734
rect 2610 2729 2656 2851
rect 2686 2733 2751 2746
rect 2510 2632 2572 2642
rect 2686 2644 2693 2733
rect 2745 2644 2751 2733
rect 2785 2720 2831 2851
rect 2958 2843 3179 2889
rect 2860 2732 2922 2742
rect 2686 2632 2751 2644
rect 2860 2640 2864 2732
rect 2918 2640 2922 2732
rect 2958 2721 3004 2843
rect 3038 2734 3103 2747
rect 2860 2630 2922 2640
rect 3038 2645 3045 2734
rect 3097 2645 3103 2734
rect 3133 2712 3179 2843
rect 3314 2851 3535 2897
rect 3214 2732 3276 2742
rect 3038 2633 3103 2645
rect 3214 2640 3218 2732
rect 3272 2640 3276 2732
rect 3314 2729 3360 2851
rect 3389 2733 3454 2746
rect 3214 2630 3276 2640
rect 3389 2644 3396 2733
rect 3448 2644 3454 2733
rect 3489 2720 3535 2851
rect 3664 2851 3885 2897
rect 3568 2734 3630 2744
rect 3389 2632 3454 2644
rect 3568 2642 3572 2734
rect 3626 2642 3630 2734
rect 3664 2729 3710 2851
rect 3568 2632 3630 2642
rect 3741 2728 3806 2741
rect 3741 2639 3748 2728
rect 3800 2639 3806 2728
rect 3839 2720 3885 2851
rect 4018 2849 4239 2895
rect 3920 2734 3982 2744
rect 3741 2627 3806 2639
rect 3920 2642 3924 2734
rect 3978 2642 3982 2734
rect 4018 2727 4064 2849
rect 4094 2728 4159 2741
rect 3920 2632 3982 2642
rect 4094 2639 4101 2728
rect 4153 2639 4159 2728
rect 4193 2718 4239 2849
rect 4367 2847 4588 2893
rect 4270 2730 4332 2740
rect 4094 2627 4159 2639
rect 4270 2638 4274 2730
rect 4328 2638 4332 2730
rect 4367 2725 4413 2847
rect 4446 2728 4511 2741
rect 4270 2628 4332 2638
rect 4446 2639 4453 2728
rect 4505 2639 4511 2728
rect 4542 2716 4588 2847
rect 4721 2851 4942 2897
rect 4624 2730 4686 2740
rect 4446 2627 4511 2639
rect 4624 2638 4628 2730
rect 4682 2638 4686 2730
rect 4721 2729 4767 2851
rect 4624 2628 4686 2638
rect 4800 2727 4865 2740
rect 4800 2638 4807 2727
rect 4859 2638 4865 2727
rect 4896 2720 4942 2851
rect 5075 2847 5296 2893
rect 4974 2732 5036 2742
rect 4800 2626 4865 2638
rect 4974 2640 4978 2732
rect 5032 2640 5036 2732
rect 5075 2725 5121 2847
rect 5149 2733 5214 2746
rect 4974 2630 5036 2640
rect 5149 2644 5156 2733
rect 5208 2644 5214 2733
rect 5250 2716 5296 2847
rect 5428 2847 5649 2893
rect 5328 2732 5390 2742
rect 5149 2632 5214 2644
rect 5328 2640 5332 2732
rect 5386 2640 5390 2732
rect 5428 2725 5474 2847
rect 5502 2728 5567 2741
rect 5328 2630 5390 2640
rect 5502 2639 5509 2728
rect 5561 2639 5567 2728
rect 5603 2716 5649 2847
rect 5679 2733 5744 2746
rect 5502 2627 5567 2639
rect 5679 2644 5686 2733
rect 5738 2644 5744 2733
rect 5679 2632 5744 2644
rect 1726 646 1772 768
rect 1901 646 1947 777
rect 1726 600 1947 646
rect 2079 644 2125 766
rect 2254 644 2300 775
rect 2079 598 2300 644
rect 2430 646 2476 768
rect 2605 646 2651 777
rect 2782 670 2828 768
rect 2957 670 3003 777
rect 2430 600 2651 646
rect 2780 600 3003 670
rect 3135 646 3181 768
rect 3310 646 3356 777
rect 3135 600 3356 646
rect 3488 646 3534 768
rect 3663 646 3709 777
rect 3488 600 3709 646
rect 3838 647 3884 769
rect 4013 647 4059 778
rect 3838 601 4059 647
rect 4193 647 4239 769
rect 4368 647 4414 778
rect 4193 601 4414 647
rect 4542 647 4588 769
rect 4717 647 4763 778
rect 4542 601 4763 647
rect 4894 646 4940 768
rect 5069 646 5115 777
rect 4894 600 5115 646
rect 5246 647 5292 769
rect 5421 647 5467 778
rect 5246 601 5467 647
rect 5599 647 5645 769
rect 5774 647 5820 778
rect 5599 601 5820 647
rect 1765 550 1895 562
rect 1765 491 1780 550
rect 1879 491 1895 550
rect 1765 44 1895 491
rect 2780 390 3000 600
rect 2780 330 2800 390
rect 2980 330 3000 390
rect 2780 310 3000 330
rect 5640 550 5780 570
rect 5640 460 5660 550
rect 5760 460 5780 550
rect 5640 90 5780 460
<< via1 >>
rect 3050 5620 3130 5680
rect 2800 5470 2852 5570
rect 3000 5470 3052 5570
rect 3190 5470 3242 5570
rect 3380 5470 3432 5570
rect 5480 5510 5532 5610
rect 5670 5510 5722 5610
rect 2720 3600 2772 3700
rect 2900 3600 2952 3700
rect 3090 3600 3142 3700
rect 3280 3600 3332 3700
rect 3470 3600 3522 3700
rect 1909 3479 1961 3540
rect 5380 3630 5432 3730
rect 5580 3630 5632 3730
rect 1810 2636 1864 2728
rect 1983 2642 2035 2731
rect 2158 2636 2212 2728
rect 2340 2644 2392 2733
rect 2514 2642 2568 2734
rect 2693 2644 2745 2733
rect 2864 2640 2918 2732
rect 3045 2645 3097 2734
rect 3218 2640 3272 2732
rect 3396 2644 3448 2733
rect 3572 2642 3626 2734
rect 3748 2639 3800 2728
rect 3924 2642 3978 2734
rect 4101 2639 4153 2728
rect 4274 2638 4328 2730
rect 4453 2639 4505 2728
rect 4628 2638 4682 2730
rect 4807 2638 4859 2727
rect 4978 2640 5032 2732
rect 5156 2644 5208 2733
rect 5332 2640 5386 2732
rect 5509 2639 5561 2728
rect 5686 2644 5738 2733
<< metal2 >>
rect 1710 5680 3140 5690
rect 1710 5620 3050 5680
rect 3130 5620 3140 5680
rect 1710 5610 3140 5620
rect 5471 5610 5731 5620
rect 2791 5570 3441 5580
rect 2791 5470 2800 5570
rect 2852 5470 3000 5570
rect 3052 5470 3190 5570
rect 3242 5470 3380 5570
rect 3432 5470 3441 5570
rect 5471 5510 5480 5610
rect 5532 5510 5670 5610
rect 5722 5510 5731 5610
rect 5471 5500 5731 5510
rect 2791 5460 2861 5470
rect 2991 5460 3061 5470
rect 3181 5460 3251 5470
rect 3371 5460 3441 5470
rect 5371 3730 5641 3740
rect 2711 3705 2781 3710
rect 2891 3705 2961 3710
rect 3081 3705 3151 3710
rect 3271 3705 3341 3710
rect 3461 3705 3531 3710
rect 2711 3700 3531 3705
rect 2711 3600 2720 3700
rect 2772 3600 2900 3700
rect 2952 3600 3090 3700
rect 3142 3600 3280 3700
rect 3332 3600 3470 3700
rect 3522 3600 3531 3700
rect 5371 3630 5380 3730
rect 5432 3630 5580 3730
rect 5632 3630 5641 3730
rect 5371 3620 5641 3630
rect 2711 3590 3531 3600
rect 2717 3587 3525 3590
rect 1278 3547 1960 3559
rect 1278 3540 1966 3547
rect 1278 3479 1909 3540
rect 1961 3479 1966 3540
rect 1278 3470 1966 3479
rect 1278 3421 1960 3470
rect 2970 2747 3160 3587
rect 5430 2747 5630 3620
rect 1817 2746 5732 2747
rect 1817 2738 5744 2746
rect 1806 2734 5744 2738
rect 1806 2733 2514 2734
rect 1806 2731 2340 2733
rect 1806 2728 1983 2731
rect 1806 2636 1810 2728
rect 1864 2642 1983 2728
rect 2035 2728 2340 2731
rect 2035 2642 2158 2728
rect 1864 2636 2158 2642
rect 2212 2644 2340 2728
rect 2392 2644 2514 2733
rect 2212 2642 2514 2644
rect 2568 2733 3045 2734
rect 2568 2644 2693 2733
rect 2745 2732 3045 2733
rect 2745 2644 2864 2732
rect 2568 2642 2864 2644
rect 2212 2640 2864 2642
rect 2918 2645 3045 2732
rect 3097 2733 3572 2734
rect 3097 2732 3396 2733
rect 3097 2645 3218 2732
rect 2918 2640 3218 2645
rect 3272 2644 3396 2732
rect 3448 2644 3572 2733
rect 3272 2642 3572 2644
rect 3626 2728 3924 2734
rect 3626 2642 3748 2728
rect 3272 2640 3748 2642
rect 2212 2639 3748 2640
rect 3800 2642 3924 2728
rect 3978 2733 5744 2734
rect 3978 2732 5156 2733
rect 3978 2730 4978 2732
rect 3978 2728 4274 2730
rect 3978 2642 4101 2728
rect 3800 2639 4101 2642
rect 4153 2639 4274 2728
rect 2212 2638 4274 2639
rect 4328 2728 4628 2730
rect 4328 2639 4453 2728
rect 4505 2639 4628 2728
rect 4328 2638 4628 2639
rect 4682 2727 4978 2730
rect 4682 2638 4807 2727
rect 4859 2640 4978 2727
rect 5032 2644 5156 2732
rect 5208 2732 5686 2733
rect 5208 2644 5332 2732
rect 5032 2640 5332 2644
rect 5386 2728 5686 2732
rect 5386 2640 5509 2728
rect 4859 2639 5509 2640
rect 5561 2644 5686 2728
rect 5738 2644 5744 2733
rect 5561 2639 5744 2644
rect 4859 2638 5744 2639
rect 2212 2636 5744 2638
rect 1806 2632 5744 2636
rect 1806 2626 1868 2632
rect 1976 2630 2041 2632
rect 2154 2626 2216 2632
rect 2860 2630 2922 2632
rect 2970 2630 3160 2632
rect 3214 2630 3276 2632
rect 3741 2627 3806 2632
rect 4094 2627 4159 2632
rect 4270 2628 4332 2632
rect 4446 2627 4511 2632
rect 4624 2628 4686 2632
rect 4800 2626 4865 2632
rect 4974 2630 5036 2632
rect 5328 2630 5390 2632
rect 5502 2627 5567 2632
use sky130_fd_pr__nfet_01v8_lvt_Q33GG7  sky130_fd_pr__nfet_01v8_lvt_Q33GG7_0
timestamp 1666367785
transform 1 0 3121 0 1 4580
box -551 -1210 551 1210
use sky130_fd_pr__nfet_01v8_lvt_TRD6KL  sky130_fd_pr__nfet_01v8_lvt_TRD6KL_0
timestamp 1666367785
transform 1 0 1931 0 1 4360
box -211 -990 211 990
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_0
timestamp 1666356932
transform 1 0 1793 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_1
timestamp 1666356932
transform 1 0 1881 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_2
timestamp 1666356932
transform 1 0 1969 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_3
timestamp 1666356932
transform 1 0 2057 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_4
timestamp 1666356932
transform 1 0 2145 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_5
timestamp 1666356932
transform 1 0 2233 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_6
timestamp 1666356932
transform 1 0 2321 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_7
timestamp 1666356932
transform 1 0 2409 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_8
timestamp 1666356932
transform 1 0 2497 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_9
timestamp 1666356932
transform 1 0 2585 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_10
timestamp 1666356932
transform 1 0 2673 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_11
timestamp 1666356932
transform 1 0 2761 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_12
timestamp 1666356932
transform 1 0 2849 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_13
timestamp 1666356932
transform 1 0 2937 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_14
timestamp 1666356932
transform 1 0 3113 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_15
timestamp 1666356932
transform 1 0 3025 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_16
timestamp 1666356932
transform 1 0 3289 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_17
timestamp 1666356932
transform 1 0 3201 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_18
timestamp 1666356932
transform 1 0 3465 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_19
timestamp 1666356932
transform 1 0 3377 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_20
timestamp 1666356932
transform 1 0 3641 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_21
timestamp 1666356932
transform 1 0 3553 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_22
timestamp 1666356932
transform 1 0 3817 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_23
timestamp 1666356932
transform 1 0 3729 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_24
timestamp 1666356932
transform 1 0 3993 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_25
timestamp 1666356932
transform 1 0 3905 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_26
timestamp 1666356932
transform 1 0 4169 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_27
timestamp 1666356932
transform 1 0 4081 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_28
timestamp 1666356932
transform 1 0 4433 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_29
timestamp 1666356932
transform 1 0 4345 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_30
timestamp 1666356932
transform 1 0 4257 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_31
timestamp 1666356932
transform 1 0 4609 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_32
timestamp 1666356932
transform 1 0 4521 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_33
timestamp 1666356932
transform 1 0 4785 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_34
timestamp 1666356932
transform 1 0 4697 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_35
timestamp 1666356932
transform 1 0 4961 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_36
timestamp 1666356932
transform 1 0 4873 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_37
timestamp 1666356932
transform 1 0 5401 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_38
timestamp 1666356932
transform 1 0 5313 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_39
timestamp 1666356932
transform 1 0 5225 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_40
timestamp 1666356932
transform 1 0 5137 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_41
timestamp 1666356932
transform 1 0 5049 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_42
timestamp 1666356932
transform 1 0 5753 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_43
timestamp 1666356932
transform 1 0 5665 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_44
timestamp 1666356932
transform 1 0 5577 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_lvt_V4M8MU  sky130_fd_pr__nfet_01v8_lvt_V4M8MU_45
timestamp 1666356932
transform 1 0 5489 0 1 1746
box -73 -1026 73 1026
use sky130_fd_pr__pfet_01v8_MGKMGH  sky130_fd_pr__pfet_01v8_MGKMGH_0
timestamp 1666367785
transform 1 0 5551 0 1 4619
box -311 -1219 311 1219
use sky130_fd_pr__res_high_po_0p35_S8HYGH  sky130_fd_pr__res_high_po_0p35_S8HYGH_0
timestamp 1666367785
transform 1 0 4481 0 1 4588
box -201 -1218 201 1218
<< labels >>
flabel metal1 1824 109 1824 109 0 FreeSans 1600 0 0 0 VRF
flabel metal2 1332 3488 1332 3490 0 FreeSans 1600 0 0 0 VB0_75
flabel metal2 3061 5510 3061 5510 0 FreeSans 1600 0 0 0 VOUT1
flabel metal2 1810 5650 1810 5650 0 FreeSans 1600 0 0 0 VB1_4
flabel metal1 5710 170 5710 170 0 FreeSans 1600 0 0 0 VSI1
flabel locali 5550 5855 5550 5855 0 FreeSans 1600 0 0 0 VDD
flabel locali 3614 127 3614 127 0 FreeSans 1600 0 0 0 VSS
flabel metal2 3030 3325 3030 3325 0 FreeSans 1600 0 0 0 VTEST1
<< end >>
