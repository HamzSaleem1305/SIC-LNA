magic
tech sky130A
magscale 1 2
timestamp 1640930396
<< metal3 >>
rect -950 3072 949 3100
rect -950 -3072 865 3072
rect 929 -3072 949 3072
rect -950 -3100 949 -3072
<< via3 >>
rect 865 -3072 929 3072
<< mimcap >>
rect -850 2960 750 3000
rect -850 -2960 -810 2960
rect 710 -2960 750 2960
rect -850 -3000 750 -2960
<< mimcapcontact >>
rect -810 -2960 710 2960
<< metal4 >>
rect 849 3072 945 3088
rect -811 2960 711 2961
rect -811 -2960 -810 2960
rect 710 -2960 711 2960
rect -811 -2961 711 -2960
rect 849 -3072 865 3072
rect 929 -3072 945 3072
rect 849 -3088 945 -3072
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -950 -3100 850 3100
string parameters w 8 l 30.0 val 494.44 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
                                                                                                                                                                   .52u l=0.06u
MI1_1-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI1_1-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI1_2-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI1_2-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI1_3-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI1_3-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND2D8 A1 A2 ZN VDD VSS
MI36 net026 A2 VSS VSS nch w=0.23u l=0.06u
MI35 ZN A1 net026 VSS nch w=0.23u l=0.06u
MI20 net032 A2 VSS VSS nch w=0.39u l=0.06u
MI17 ZN A1 net032 VSS nch w=0.39u l=0.06u
MI21 net031 A2 VSS VSS nch w=0.39u l=0.06u
MI23 ZN A1 net050 VSS nch w=0.39u l=0.06u
MI22 ZN A1 net031 VSS nch w=0.39u l=0.06u
MI26 ZN A1 net053 VSS nch w=0.39u l=0.06u
MI19 ZN A1 net071 VSS nch w=0.39u l=0.06u
MI24 net050 A2 VSS VSS nch w=0.39u l=0.06u
MI25 net053 A2 VSS VSS nch w=0.39u l=0.06u
MI27 ZN A1 net059 VSS nch w=0.39u l=0.06u
MI28 net059 A2 VSS VSS nch w=0.39u l=0.06u
MI29 net062 A2 VSS VSS nch w=0.23u l=0.06u
MI18 net071 A2 VSS VSS nch w=0.39u l=0.06u
MI30 ZN A1 net062 VSS nch w=0.23u l=0.06u
M_u2_0 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_1 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_2 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_3 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_4 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_5 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_6 ZN A2 VDD VDD pch w=0.52u l=0.06u
M_u2_7 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI6_0 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_2 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_3 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_4 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_5 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_6 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI6_7 ZN A1 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND3D0 A1 A2 A3 ZN VDD VSS
MI0-M_u4 ZN A1 XI0-net10 VSS nch w=0.195u l=0.06u
MI0-M_u5 XI0-net10 A2 XI0-net13 VSS nch w=0.195u l=0.06u
MI0-M_u6 XI0-net13 A3 VSS VSS nch w=0.195u l=0.06u
MI0-M_u3 ZN A3 VDD VDD pch w=0.26u l=0.06u
MI0-M_u1 ZN A1 VDD VDD pch w=0.26u l=0.06u
MI0-M_u2 ZN A2 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt ND3D1 A1 A2 A3 ZN VDD VSS
MI1-M_u4 ZN A1 XI1-net10 VSS nch w=0.39u l=0.06u
MI1-M_u5 XI1-net10 A2 XI1-net13 VSS nch w=0.39u l=0.06u
MI1-M_u6 XI1-net13 A3 VSS VSS nch w=0.39u l=0.06u
MI1-M_u3 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI1-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI1-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND3D2 A1 A2 A3 ZN VDD VSS
MI0_0-M_u4 ZN A1 XI0_0-net10 VSS nch w=0.39u l=0.06u
MI0_0-M_u5 XI0_0-net10 A2 XI0_0-net13 VSS nch w=0.39u l=0.06u
MI0_0-M_u6 XI0_0-net13 A3 VSS VSS nch w=0.39u l=0.06u
MI0_1-M_u4 ZN A1 XI0_1-net10 VSS nch w=0.39u l=0.06u
MI0_1-M_u5 XI0_1-net10 A2 XI0_1-net13 VSS nch w=0.39u l=0.06u
MI0_1-M_u6 XI0_1-net13 A3 VSS VSS nch w=0.39u l=0.06u
MI0_0-M_u3 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI0_0-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI0_0-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI0_1-M_u3 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI0_1-M_u1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI0_1-M_u2 ZN A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND3D3 A1 A2 A3 ZN VDD VSS
MI0_0-M_u4 ZN A1 XI0_0-net10 VSS nch w=0.39u l=0.06u
MI0_0-M_u5 XI0_0-net10 A2 XI0_0-timestamp 1640952342
version 8.3
tech sky130A
style ngspice()
scale 1000 1 500000
resistclasses 4400000 2200000 1700000 3050000 120000 197000 114000 191000 120000 197000 114000 191000 48200 319800 2000000 48200 48200 12200 125 125 47 47 29 5
parameters sky130_fd_pr__cap_mim_m3_1 w=w l=l
node "c1_n3050_n1000#" 0 0 -3050 -1000 mim 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 11382084 15688 0 0 0 0
node "m3_n3150_n1100#" 1 7641.93 -3150 -1100 m3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13857800 16998 208896 4544 0 0 0 0
substrate "VSUBS" 0 0 -1073741817 -1073741817 space 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
cap "m3_n3150_n1100#" "c1_n3050_n1000#" 30404.8
device csubckt sky130_fd_pr__cap_mim_m3_1 -3050 -1000 -3049 -999 w=6000 l=2000 "None" "c1_n3050_n1000#" 15680 0 "m3_n3150_n1100#" 2840 0
                                                                                          6u
MI12_1 ZN A1 net24<1> VSS nch w=0.39u l=0.06u
MI12_2 ZN A1 net24<2> VSS nch w=0.39u l=0.06u
MI12_3 ZN A1 net24<3> VSS nch w=0.39u l=0.06u
MI5_0 net21<0> A3 VSS VSS nch w=0.39u l=0.06u
MI5_1 net21<1> A3 VSS VSS nch w=0.39u l=0.06u
MI5_2 net21<2> A3 VSS VSS nch w=0.39u l=0.06u
MI5_3 net21<3> A3 VSS VSS nch w=0.39u l=0.06u
MI2_0 net24<0> A2 net21<0> VSS nch w=0.39u l=0.06u
MI2_1 net24<1> A2 net21<1> VSS nch w=0.39u l=0.06u
MI2_2 net24<2> A2 net21<2> VSS nch w=0.39u l=0.06u
MI2_3 net24<3> A2 net21<3> VSS nch w=0.39u l=0.06u
.ends
.subckt ND3D8 A1 A2 A3 ZN VDD VSS
MI0-M_u4 ZN A1 XI0-net10 VSS nch w=3.12u l=0.06u
MI0-M_u5 XI0-net10 A2 XI0-net13 VSS nch w=3.12u l=0.06u
MI0-M_u6 XI0-net13 A3 VSS VSS nch w=3.12u l=0.06u
MI0-M_u3 ZN A3 VDD VDD pch w=4.16u l=0.06u
MI0-M_u1 ZN A1 VDD VDD pch w=4.16u l=0.06u
MI0-M_u2 ZN A2 VDD VDD pch w=4.16u l=0.06u
.ends
.subckt ND4D0 A1 A2 A3 A4 ZN VDD VSS
MI19 p2 A4 VSS VSS nch w=0.195u l=0.06u
MI17 p0 A2 p1 VSS nch w=0.195u l=0.06u
MI18 p1 A3 p2 VSS nch w=0.195u l=0.06u
MU53 ZN A1 p0 VSS nch w=0.195u l=0.06u
MI14 ZN A3 VDD VDD pch w=0.26u l=0.06u
MI15 ZN A2 VDD VDD pch w=0.26u l=0.06u
MI16 ZN A1 VDD VDD pch w=0.26u l=0.06u
MI9 ZN A4 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt ND4D1 A1 A2 A3 A4 ZN VDD VSS
MI5 p2 A4 VSS VSS nch w=0.39u l=0.06u
MI3 p0 A2 p1 VSS nch w=0.39u l=0.06u
MI4 p1 A3 p2 VSS nch w=0.39u l=0.06u
MU53 ZN A1 p0 VSS nch w=0.39u l=0.06u
MI7 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI2 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI1 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI0 ZN A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND4D2 A1 A2 A3 A4 ZN VDD VSS
MI12_0 p2 A4 VSS VSS nch w=0.39u l=0.06u
MI12_1 p2 A4 VSS VSS nch w=0.39u l=0.06u
MI9_0 p0 A2 p1 VSS nch w=0.39u l=0.06u
MI9_1 p0 A2 p1 VSS nch w=0.39u l=0.06u
MI11_0 p1 A3 p2 VSS nch w=0.39u l=0.06u
MI11_1 p1 A3 p2 VSS nch w=0.39u l=0.06u
MU53_0 ZN A1 p0 VSS nch w=0.39u l=0.06u
MU53_1 ZN A1 p0 VSS nch w=0.39u l=0.06u
MI8_0 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI8_1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI2_0 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI2_1 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI6_0 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI6_1 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI7_0 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI7_1 ZN A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND4D3 A1 A2 A3 A4 ZN VDD VSS
MI28 net026 A3 net023 VSS nch w=1.17u l=0.06u
MI29 net023 A4 VSS VSS nch w=1.17u l=0.06u
MI27 net029 A2 net026 VSS nch w=1.17u l=0.06u
MU53 ZN A1 net029 VSS nch w=1.17u l=0.06u
MI8_0 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI8_1 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI8_2 ZN A1 VDD VDD pch w=0.52u l=0.06u
MI2_0 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI2_1 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI2_2 ZN A4 VDD VDD pch w=0.52u l=0.06u
MI6_0 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI6_1 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI6_2 ZN A3 VDD VDD pch w=0.52u l=0.06u
MI7_0 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI7_1 ZN A2 VDD VDD pch w=0.52u l=0.06u
MI7_2 ZN A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ND4D4 A1 A2 A3 A4 ZN VDD VSS
MU3-M_u5 ZN A1 XU3-net23 VSS nch w=1.56u l=0.06u
MU3-MI0 XU3-net23 A2 XU3-net26 VSS nch w=1.5timestamp 1640943879
version 8.3
tech sky130A
style ngspice()
scale 1000 1 500000
resistclasses 4400000 2200000 1700000 3050000 120000 197000 114000 191000 120000 197000 114000 191000 48200 319800 2000000 48200 48200 12200 125 125 47 47 29 5
use CurrentMirror_layout CurrentMirror_layout_0 1 0 634 0 1 -2505
use DiffPair_layout DiffPair_layout_0 1 0 462 0 1 701
use sky130_fd_pr__cap_mim_m3_1_TQVBRR sky130_fd_pr__cap_mim_m3_1_TQVBRR_0 1 0 8075 0 1 -2427
use PMOS2 PMOS2_0 1 0 4139 0 1 1699
use PMOS_Load PMOS_Load_0 1 0 490 0 1 3052
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1 1 0 8671 0 1 6190
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 -1 0 2036 0 1 6190
node "IBIAS" 2 6962.43 -9176 -858 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 6391705 20712 0 0 0 0 0 0 0 0
node "m2_1498_1216#" 1 1227.97 1498 1216 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56184 1370 567250 5038 0 0 0 0 0 0
node "m2_864_n933#" 1 1227.97 864 -933 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56184 1370 567250 5038 0 0 0 0 0 0
node "VO" 3 17392 2108 -2389 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 8439882 25440 1307826 6480 28921181 37724 0 0 0 0
node "m2_3531_794#" 1 1429.39 3531 794 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13770 664 586460 5442 0 0 0 0 0 0
node "m2_530_794#" 1 1398.62 530 794 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13770 664 586460 5442 0 0 0 0 0 0
node "m2_2582_1554#" 2 1436.04 2582 1554 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 17800 756 359568 5712 0 0 0 0 0 0
node "m2_1003_1555#" 2 1407.26 1003 1555 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 17800 756 359568 5712 0 0 0 0 0 0
node "VN" 2 7814.79 -1045 241 m1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 675091 4720 6308515 19544 0 0 0 0 0 0 0 0
node "VP" 3 7814.27 -584 1496 m1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 391624 4952 6308515 19544 0 0 0 0 0 0 0 0
node "m1_5404_4055#" 2 7061.38 5404 4055 m1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 36720 772 180700 3310 4955840 15936 10899636 13990 0 0 0 0
node "VSS" 81 122646 107 -163 li 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 7756104 16428 794626 4030 112073122 106086 110747267 125354 15446591 30328 0 0 0 0
node "VDD" 214 94485.9 536 4549 li 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 7778407 24572 5663175 20848 88011407 88620 64944036 92864 31012240 26472 0 0 0 0
node "w_5404_4055#" 2160 110.16 5404 4055 nw 0 0 0 0 36720 772 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
substrate "VSUBS" 0 0 -1073741817 -1073741817 space 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
cap "VDD" "VSS" 31319
cap "m2_864_n933#" "m2_530_794#" 230.436
cap "m1_5404_4055#" "VO" 4792.46
cap "VDD" "IBIAS" 3797.94
cap "VSS" "IBIAS" 4767
cap "m2_1498_1216#" "VSS" 363.377
cap "m2_1003_1555#" "VDD" 15.4514
cap "VDD" "VP" 3797.94
cap "VDD" "VN" 3797.94
cap "VP" "VSS" 4767
cap "VN" "VSS" 4767
cap "w_5404_4055#" "m1_5404_4055#" 23.868
cap "VDD" "VO" 12104.1
cap "VO" "VSS" 15801.2
cap "m2_864_n933#" "VSS" 363.377
cap "VDD" "m1_5404_4055#" 2320.81
cap "m2_1003_1555#" "VP" 78.232
cap "VDD" "m2_2582_1554#" 15.614
cap "m2_1498_1216#" "m2_864_n933#" 374.207
cap "m2_1003_1555#" "m2_864_n933#" 43.3298
cap "m2_1003_1555#" "m2_530_794#" 368.324
cap "m2_530_794#" "VP" 112.136
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" 51.3197
cap "CurrentMirror_layout_0/D3" "CurrentMirror_layout_0/S" 698.143
cap "CurrentMirror_layout_0/D1" "CurrentMirror_layout_0/S" 3.22744
cap "CurrentMirror_layout_0/D3" "CurrentMirror_layout_0/D1" 690.375
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 1610.1
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 262.005
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "VO" -246.231
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 2653.96
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -527.1
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "VO" -575.025
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "VO" 2653.96
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -101.02
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -234.29
cap "CurrentMirror_layout_0/S" "CurrentMirror_layout_0/D1" 284.196
cap "CurrentMirror_layout_0/S" "CurrentMirror_layout_0/D2" 704.237
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_7/a_50_n1050#" "CurrentMirror_layout_0/D2" 2.84217e-14
cap "CurrentMirror_layout_0/D1" "CurrentMirror_layout_0/D2" 2100.43
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_0/a_n108_n1050#" "CurrentMirror_layout_0/D2" 1.13687e-13
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_3/a_50_n1050#" "CurrentMirror_layout_0/D2" 2.27374e-13
cap "CurrentMirror_layout_0/S" "VO" 77.5641
cap "CurrentMirror_layout_0/S" "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_5/a_n50_n1076#" 3.22744
cap "CurrentMirror_layout_0/S" "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_9/a_50_n1050#" 87.2639
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_5/a_n50_n1076#" "CurrentMirror_layout_0/D2" -82.205
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_9/a_50_n1050#" "CurrentMirror_layout_0/D2" -2.84217e-14
cap "m1_5404_4055#" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 190.612
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/w_n389_n527#" 322.73
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 2.13163e-14
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -98.6
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/G1" 66.7336
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 187.705
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -80.8235
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/w_n389_n527#" 401.3
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 493.62
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 1017.21
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_6/a_n50_n526#" 221.055
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_2/a_n50_n526#" 221.055
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 4.54747e-13
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_18/a_n50_n526#" 185.639
cap "m1_5404_4055#" "PMOS2_0/S" 38.8284
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/D1" 51.65
cap "m1_5404_4055#" "DiffPair_layout_0/w_n389_n527#" 613.17
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 222.724
cap "PMOS2_0/S" "m1_5404_4055#" 5.3352
cap "PMOS2_0/S" "VO" 18.9696
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -315.819
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/G2" 322.73
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -15.6202
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 90.195
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -96.8202
cap "PMOS_Load_0/S" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 3.06
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 7.8859
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 216.993
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 111.527
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" -23.985
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_3/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 42.74
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 36.485
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 214.483
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -72.9359
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_7/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 42.74
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 252.378
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_3/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 52.3
cap "PMOS_Load_0/S" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 3.366
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 98.1339
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 57.2455
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 89.92
cap "PMOS_Load_0/S" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 2.958
cap "DiffPair_layout_0/S" "DiffPair_layout_0/D1" -132.44
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/D2" 216.912
cap "PMOS_Load_0/S" "DiffPair_layout_0/D2" 3.366
cap "DiffPair_layout_0/S" "DiffPair_layout_0/D2" 112.045
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/D1" -51
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/D2" -198.66
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/D2" 252.378
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_19/a_n50_n526#" "DiffPair_layout_0/D1" 16.85
cap "DiffPair_layout_0/D1" "PMOS_Load_0/S" 6.018
cap "PMOS_Load_0/S" "m1_5404_4055#" 58.641
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 472.795
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/D1" 315.028
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/w_n389_n527#" 281.355
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/D2" 223.993
cap "DiffPair_layout_0/w_n389_n527#" "m1_5404_4055#" 648.543
cap "PMOS2_0/S" "m1_5404_4055#" 7.56
cap "PMOS2_0/G" "PMOS2_0/D" 897.876
cap "PMOS2_0/S" "PMOS2_0/D" 622.285
cap "PMOS2_0/S" "VO" -203.047
cap "PMOS_Load_0/D1" "PMOS_Load_0/S" -99.4994
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" 1139.21
cap "PMOS_Load_0/S" "PMOS_Load_0/D1" 126.929
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 786.318
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" 967.005
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 200.884
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" "PMOS_Load_0/D2" 585.435
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" 172.201
cap "PMOS_Load_0/D1" "PMOS_Load_0/D1" -73.68
cap "PMOS_Load_0/D2" "PMOS_Load_0/D1" -1.44
cap "PMOS_Load_0/S" "PMOS_Load_0/D1" 337.38
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 384.612
cap "PMOS2_0/G" "PMOS2_0/S" 118.104
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n108_n600#" "PMOS_Load_0/S" 8.04255
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 7.73381
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 24.35
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/S" 142.558
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" "PMOS_Load_0/S" 18.7864
cap "PMOS_Load_0/D2" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_7/a_50_n600#" 5.68434e-14
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_7/a_50_n600#" 8.80851
cap "PMOS_Load_0/D2" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n108_n600#" -82.205
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 413.144
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1564.78
cap "PMOS_Load_0/D2" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_3/a_50_n600#" -2.27374e-13
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_3/a_50_n600#" "PMOS_Load_0/S" 8.80851
cap "PMOS_Load_0/D2" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" 268.73
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" "PMOS_Load_0/S" 611.65
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 131.82
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_n50_n626#" "PMOS_Load_0/S" 611.65
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1384.48
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 261.66
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_n50_n626#" "PMOS_Load_0/D2" 268.73
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_16/a_n108_n600#" 8.80851
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" "PMOS_Load_0/S" 39.2553
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 49.32
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_12/a_n108_n600#" 8.80851
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" "PMOS_Load_0/D2" 155.002
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 56.54
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -12.32
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_19/a_50_n600#" 8.80851
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_15/a_n50_n626#" 215.825
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1384.48
cap "PMOS2_0/S" "PMOS2_0/G" 175.002
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS2_0/S" -206.885
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 57.5463
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "PMOS2_0/S" -14.85
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "PMOS2_0/S" 1261.4
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "PMOS2_0/S" 49.32
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "PMOS2_0/S" 1384.48
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "PMOS2_0/S" 49.32
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1384.48
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 63.55
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1204.02
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" -1352.34
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 117.549
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 154
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 386.26
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "VDD" -1378.37
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 4067.93
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 3985.43
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 3985.43
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1486.5
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 253.499
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 253.499
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" -870.93
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 263.284
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 2470.58
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "VDD" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 4239.25
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "VDD" -1240.4
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 453.67
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 518.775
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 70.11
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 386.8
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1645.15
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 2187.5
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 2443
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 2538.14
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 854.147
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 1561.69
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 92.9015
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 2443
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 2443
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 2241.96
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1111.78
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" -70.3871
merge "PMOS_Load_0/D1" "DiffPair_layout_0/D1" -1862.94 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -138970 -1328 -373736 -3878 0 0 0 0 0 0
merge "DiffPair_layout_0/D1" "m2_3531_794#"
merge "m2_3531_794#" "m2_530_794#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/VSUBS" -11197.3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -5394990 -20718 0 0 0 0 0 0 -777170 -11492 0 0 0 0
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/VSUBS" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/VSUBS"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/VSUBS" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/VSUBS"
merge "PMOS_Load_0/VSUBS" "PMOS2_0/VSUBS"
merge "PMOS2_0/VSUBS" "DiffPair_layout_0/w_n389_n527#"
merge "DiffPair_layout_0/w_n389_n527#" "CurrentMirror_layout_0/S"
merge "CurrentMirror_layout_0/S" "VSS"
merge "VSS" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/VSUBS"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/VSUBS" "VSUBS"
merge "PMOS2_0/G" "PMOS_Load_0/D2" -4296.62 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 3335 -472 -935032 -2260 48840 -2230 0 0 0 0 0 0
merge "PMOS_Load_0/D2" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "m1_5404_4055#"
merge "m1_5404_4055#" "DiffPair_layout_0/D2"
merge "DiffPair_layout_0/D2" "m2_2582_1554#"
merge "m2_2582_1554#" "m2_1003_1555#"
merge "DiffPair_layout_0/S" "CurrentMirror_layout_0/D2" -2812.1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -24247 -2740 -306139 -6596 0 0 0 0 0 0
merge "CurrentMirror_layout_0/D2" "m2_1498_1216#"
merge "m2_1498_1216#" "m2_864_n933#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -38606 0 0 0 0 -26690 -772 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -605657 -26722 1466048 -14587 -26748840 -32187 -2287682 -27214 -21157388 -26923 0 0 0 0
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS_Load_0/S"
merge "PMOS_Load_0/S" "w_5404_4055#"
merge "w_5404_4055#" "PMOS2_0/S"
merge "PMOS2_0/S" "VDD"
merge "PMOS2_0/D" "CurrentMirror_layout_0/D3" -11174.6 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -4857782 -20481 -3468453 -7600 -913924 -20467 0 0 0 0
merge "CurrentMirror_layout_0/D3" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "VO"
merge "DiffPair_layout_0/G1" "VN" 170.229 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 161075 -328 167475 0 0 0 0 0 0 0 0 0
merge "DiffPair_layout_0/G2" "VP" -475.348 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -26880 -1166 0 0 0 0 0 0 0 0 0 0
merge "CurrentMirror_layout_0/D1" "IBIAS" -476.836 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -452007 -342 0 0 0 0 0 0 0 0
                                                                                                                                                                                                                                                                                                                                                                                                       et36 A1 net27 VSS nch w=0.39u l=0.06u
MU25 net39 C1 VSS VSS nch w=0.39u l=0.06u
MI19_0-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI19_1-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI8 net36 C2 net46 VDD pch w=0.52u l=0.06u
MI2 net46 C1 VDD VDD pch w=0.52u l=0.06u
MI13 net36 A1 net34 VDD pch w=0.52u l=0.06u
MI12 net34 A2 VDD VDD pch w=0.52u l=0.06u
MI9 net36 B2 net37 VDD pch w=0.52u l=0.06u
MI11 net37 B1 VDD VDD pch w=0.52u l=0.06u
MI19_0-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
MI19_1-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt OA222D4 A1 A2 B1 B2 C1 C2 Z VDD VSS
MI34 net36 A2 net27 VSS nch w=0.78u l=0.06u
MI30 net39 C2 VSS VSS nch w=0.78u l=0.06u
MI31 net27 B1 net39 VSS nch w=0.78u l=0.06u
MI32 net27 B2 net39 VSS nch w=0.78u l=0.06u
MI33 net36 A1 net27 VSS nch w=0.78u l=0.06u
MI29 net39 C1 VSS VSS nch w=0.78u l=0.06u
MI19_0-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI19_1-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI19_2-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI19_3-M_u2 Z net36 VSS VSS nch w=0.39u l=0.06u
MI23_0 net57<0> C1 VDD VDD pch w=0.52u l=0.06u
MI23_1 net57<1> C1 VDD VDD pch w=0.52u l=0.06u
MI24_0 net36 C2 net57<0> VDD pch w=0.52u l=0.06u
MI24_1 net36 C2 net57<1> VDD pch w=0.52u l=0.06u
MI20_0 net36 A1 net69<0> VDD pch w=0.52u l=0.06u
MI20_1 net36 A1 net69<1> VDD pch w=0.52u l=0.06u
MI12_0 net69<0> A2 VDD VDD pch w=0.52u l=0.06u
MI12_1 net69<1> A2 VDD VDD pch w=0.52u l=0.06u
MI21_0 net36 B2 net66<0> VDD pch w=0.52u l=0.06u
MI21_1 net36 B2 net66<1> VDD pch w=0.52u l=0.06u
MI22_0 net66<0> B1 VDD VDD pch w=0.52u l=0.06u
MI22_1 net66<1> B1 VDD VDD pch w=0.52u l=0.06u
MI19_0-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
MI19_1-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
MI19_2-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
MI19_3-M_u3 Z net36 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt OA22D0 A1 A2 B1 B2 Z VDD VSS
M_u4 net29 B2 VSS VSS nch w=0.195u l=0.06u
MI19 net30 A2 net29 VSS nch w=0.195u l=0.06u
MI20 net30 A1 net29 VSS nch w=0.195u l=0.06u
MI18 net29 B1 VSS VSS nch w=0.195u l=0.06u
MU1-M_u2 Z net30 VSS VSS nch w=0.195u l=0.06u
MU24 net25 B2 VDD VDD pch w=0.26u l=0.06u
MI16 net22 A2 VDD VDD pch w=0.26u l=0.06u
MI15 net30 B1 net25 VDD pch w=0.26u l=0.06u
MI17 net30 A1 net22 VDD pch w=0.26u l=0.06u
MU1-M_u3 Z net30 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt OA22D1 A1 A2 B1 B2 Z VDD VSS
M_u4 net29 B2 VSS VSS nch w=0.39u l=0.06u
MI13 net30 A2 net29 VSS nch w=0.39u l=0.06u
MI14 net30 A1 net29 VSS nch w=0.39u l=0.06u
MI12 net29 B1 VSS VSS nch w=0.39u l=0.06u
MU1-M_u2 Z net30 VSS VSS nch w=0.39u l=0.06u
MU24 net25 B2 VDD VDD pch w=0.52u l=0.06u
MI11 net22 A2 VDD VDD pch w=0.52u l=0.06u
MI8 net30 B1 net25 VDD pch w=0.52u l=0.06u
MI9 net30 A1 net22 VDD pch w=0.52u l=0.06u
MU1-M_u3 Z net30 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt OA22D2 A1 A2 B1 B2 Z VDD VSS
M_u4 net29 B2 VSS VSS nch w=0.39u l=0.06u
MI13 net30 A2 net29 VSS nch w=0.39u l=0.06u
MI14 net30 A1 net29 VSS nch w=0.39u l=0.06u
MI12 net29 B1 VSS VSS nch w=0.39u l=0.06u
MU1_0-M_u2 Z net30 VSS VSS nch w=0.39u l=0.06u
MU1_1-M_u2 Z net30 VSS VSS nch w=0.39u l=0.06u
MU24 net2* NGSPICE file created from OpampM.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_RC9KLY a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS
X0 a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=500000u
.ends

.subckt CurrentMirror_layout D3 D2 D1 S
Xsky130_fd_pr__nfet_01v8_RC9KLY_1 D2 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_3 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_2 S D1 D2 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_4 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_5 D1 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_6 S D1 D1 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_7 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_8 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_9 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_0 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
.ends

.subckt sky130_fd_pr__nfet_01v8_6YBK2C a_50_n500# a_n50_n526# a_n108_n500# VSUBS
X0 a_50_n500# a_n50_n526# a_n108_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt DiffPair_layout D2 D1 G2 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
Xsky130_fd_pr__nfet_01v8_6YBK2C_10 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_11 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_13 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_12 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_14 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_15 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_16 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_17 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_18 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_19 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_0 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_2 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_1 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_3 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_4 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_5 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_6 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_7 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_8 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_9 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_EEU9S7 w_n144_n662# a_50_n600# a_n50_n626#
+ a_n108_n600# VSUBS
X0 a_50_n600# a_n50_n626# a_n108_n600# w_n144_n662# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
.ends

.subckt PMOS_Load D2 D1 S VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_0 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_1 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_10 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_2 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_11 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_3 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_12 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_4 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_13 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_5 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_14 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_7 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_6 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_15 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_8 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_16 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_9 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_17 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_19 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_18 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TQVBRR m3_n2550_n2500# c1_n2450_n2400# VSUBS
X0 c1_n2450_n2400# m3_n2550_n2500# sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.4e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_N3PKNJ c1_n3050_n1000# m3_n3150_n1100# VSUBS
X0 c1_n3050_n1000# m3_n3150_n1100# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_WFBLZ7 a_50_n1420# a_n50_n1446# w_n144_n1482# a_n108_n1420#
+ VSUBS
X0 a_50_n1420# a_n50_n1446# a_n108_n1420# w_n144_n1482# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.42e+07u l=500000u
.ends

.subckt PMOS2 G D S VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_19 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_0 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_1 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_2 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_3 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_5 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_4 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_6 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_7 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_8 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_9 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_20 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_21 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_10 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_22 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_11 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_23 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_12 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_24 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_13 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_14 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_15 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_16 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_17 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_18 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
.ends


* Top level circuit OpampM

XCurrentMirror_layout_0 VO DiffPair_layout_0/S IBIAS VSS CurrentMirror_layout
XDiffPair_layout_0 PMOS2_0/G PMOS_Load_0/D1 VP VN DiffPair_layout_0/S VSS DiffPair_layout
XPMOS_Load_0 PMOS2_0/G PMOS_Load_0/D1 VDD VSS PMOS_Load
Xsky130_fd_pr__cap_mim_m3_1_TQVBRR_0 VO PMOS2_0/G VSS sky130_fd_pr__cap_mim_m3_1_TQVBRR
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 VDD VSS VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_1 VDD VSS VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
XPMOS2_0 PMOS2_0/G VO VDD VSS PMOS2
.end

                                                                                                                                                                                        SS nch w=0.78u l=0.06u
MI22 net15 B3 VSS VSS nch w=0.78u l=0.06u
MI21 net31 A1 net15 VSS nch w=0.78u l=0.06u
MU1_0-M_u2 Z net31 VSS VSS nch w=0.39u l=0.06u
MU1_1-M_u2 Z net31 VSS VSS nch w=0.39u l=0.06u
MU1_2-M_u2 Z net31 VSS VSS nch w=0.39u l=0.06u
MU1_3-M_u2 Z net31 VSS VSS nch w=0.39u l=0.06u
MI13_0-MI12 net31 B3 XI13_0-net11 VDD pch w=0.52u l=0.06u
MI13_0-MI13 XI13_0-net11 B2 XI13_0-net18 VDD pch w=0.52u l=0.06u
MI13_0-MI15 XI13_0-net18 B1 VDD VDD pch w=0.52u l=0.06u
MI13_1-MI12 net31 B3 XI13_1-net11 VDD pch w=0.52u l=0.06u
MI13_1-MI13 XI13_1-net11 B2 XI13_1-net18 VDD pch w=0.52u l=0.06u
MI13_1-MI15 XI13_1-net18 B1 VDD VDD pch w=0.52u l=0.06u
MI19_0-MI12 net31 A3 XI19_0-net11 VDD pch w=0.52u l=0.06u
MI19_0-MI13 XI19_0-net11 A2 XI19_0-net18 VDD pch w=0.52u l=0.06u
MI19_0-MI15 XI19_0-net18 A1 VDD VDD pch w=0.52u l=0.06u
MI19_1-MI12 net31 A3 XI19_1-net11 VDD pch w=0.52u l=0.06u
MI19_1-MI13 XI19_1-net11 A2 XI19_1-net18 VDD pch w=0.52u l=0.06u
MI19_1-MI15 XI19_1-net18 A1 VDD VDD pch w=0.52u l=0.06u
MU1_0-M_u3 Z net31 VDD VDD pch w=0.52u l=0.06u
MU1_1-M_u3 Z net31 VDD VDD pch w=0.52u l=0.06u
MU1_2-M_u3 Z net31 VDD VDD pch w=0.52u l=0.06u
MU1_3-M_u3 Z net31 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt OAI211D0 A1 A2 B C ZN VDD VSS
MI8 net36 B net24 VSS nch w=0.195u l=0.06u
MI9 net24 C VSS VSS nch w=0.195u l=0.06u
M_u2 ZN A1 net36 VSS nch w=0.195u l=0.06u
MI7 ZN A2 net36 VSS nch w=0.195u l=0.06u
MI6 ZN A2 net35 VDD pch w=0.26u l=0.06u
MI5 net35 A1 VDD VDD pch w=0.26u l=0.06u
MI4 ZN C VDD VDD pch w=0.26u l=0.06u
M_u12 ZN B VDD VDD pch w=0.26u l=0.06u
.ends
.subckt OAI211D1 A1 A2 B C ZN VDD VSS
MI2 net36 B net24 VSS nch w=0.39u l=0.06u
MI3 net24 C VSS VSS nch w=0.39u l=0.06u
M_u2 ZN A1 net36 VSS nch w=0.39u l=0.06u
M_u3 ZN A2 net36 VSS nch w=0.39u l=0.06u
MI1 ZN A2 net35 VDD pch w=0.52u l=0.06u
MI0 net35 A1 VDD VDD pch w=0.52u l=0.06u
M_u11 ZN C VDD VDD pch w=0.52u l=0.06u
M_u12 ZN B VDD VDD pch w=0.52u l=0.06u
.ends
.subckt OAI211D2 A1 A2 B C ZN VDD VSS
MI8_0 net36 B net25<0> VSS nch w=0.39u l=0.06u
MI8_1 net36 B net25<1> VSS nch w=0.39u l=0.06u
MI11_0 net25<0> C VSS VSS nch w=0.39u l=0.06u
MI11_1 net25<1> C VSS VSS nch w=0.39u l=0.06u
M_u2 ZN A1 net36 VSS nch w=0.78u l=0.06u
MI13 ZN A2 net36 VSS nch w=0.78u l=0.06u
MI12_0 ZN A2 net38<0> VDD pch w=0.52u l=0.06u
MI12_1 ZN A2 net38<1> VDD pch w=0.52u l=0.06u
MI5_0 net38<0> A1 VDD VDD pch w=0.52u l=0.06u
MI5_1 net38<1> A1 VDD VDD pch w=0.52u l=0.06u
MI4 ZN C VDD VDD pch w=1.04u l=0.06u
M_u12 ZN B VDD VDD pch w=1.04u l=0.06u
.ends
.subckt OAI211D4 A1 A2 B C ZN VDD VSS
MI21 net33 B net25 VSS nch w=1.56u l=0.06u
MI22 net25 C VSS VSS nch w=1.56u l=0.06u
M_u2 ZN A1 net33 VSS nch w=1.56u l=0.06u
MI20 ZN A2 net33 VSS nch w=1.56u l=0.06u
MI19 ZN A2 net44 VDD pch w=2.08u l=0.06u
MI18 net44 A1 VDD VDD pch w=2.08u l=0.06u
MI17 ZN C VDD VDD pch w=2.08u l=0.06u
MI16 ZN B VDD VDD pch w=2.08u l=0.06u
.ends
.subckt OAI21D0 A1 A2 B ZN VDD VSS
M_u2 ZN A1 net15 VSS nch w=0.195u l=0.06u
M_u3 ZN A2 net15 VSS nch w=0.195u l=0.06u
M_u4 net15 B VSS VSS nch w=0.195u l=0.06u
M_u9 ZN B VDD VDD pch w=0.26timestamp 1640952342
version 8.3
tech sky130A
style ngspice()
scale 1000 1 500000
resistclasses 4400000 2200000 1700000 3050000 120000 197000 114000 191000 120000 197000 114000 191000 48200 319800 2000000 48200 48200 12200 125 125 47 47 29 5
use PMOS_Load PMOS_Load_0 1 0 490 0 1 3052
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 -1 0 2036 0 1 6190
use sky130_fd_pr__cap_mim_m3_1_N3PKNJ sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1 1 0 8671 0 1 6190
use PMOS2 PMOS2_0 1 0 4139 0 1 1699
use sky130_fd_pr__cap_mim_m3_1_TQVBRR sky130_fd_pr__cap_mim_m3_1_TQVBRR_0 1 0 8075 0 1 -2427
use DiffPair_layout DiffPair_layout_0 1 0 462 0 1 701
use CurrentMirror_layout CurrentMirror_layout_0 1 0 634 0 1 -2505
port "IBIAS" 6 -8852 -591 -8852 -591 m2
port "VO" 3 19494 -84 19494 -84 m4
port "VN" 5 -8791 531 -8791 531 m2
port "VP" 4 -8568 1903 -8568 1903 m2
port "VSS" 1 5268 10390 5268 10390 m2
port "VDD" 2 5485 7900 5485 7900 v2
node "IBIAS" 2 6962.43 -8852 -591 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 6391705 20712 0 0 0 0 0 0 0 0
node "m2_1498_1216#" 1 1227.97 1498 1216 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56184 1370 567250 5038 0 0 0 0 0 0
node "m2_864_n933#" 1 1227.97 864 -933 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 56184 1370 567250 5038 0 0 0 0 0 0
node "VO" 3 17341.2 19494 -84 m4 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 8439882 25440 1307826 6480 27914951 37354 0 0 0 0
node "m2_3531_794#" 1 1429.39 3531 794 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13770 664 586460 5442 0 0 0 0 0 0
node "m2_530_794#" 1 1398.62 530 794 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13770 664 586460 5442 0 0 0 0 0 0
node "m2_2582_1554#" 2 1436.04 2582 1554 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 17800 756 359568 5712 0 0 0 0 0 0
node "m2_1003_1555#" 2 1407.26 1003 1555 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 17800 756 359568 5712 0 0 0 0 0 0
node "VN" 2 7814.79 -8791 531 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 675091 4720 6308515 19544 0 0 0 0 0 0 0 0
node "VP" 3 7814.27 -8568 1903 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 391624 4952 6308515 19544 0 0 0 0 0 0 0 0
node "m1_5404_4055#" 2 7061.38 5404 4055 m1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 36720 772 180700 3310 4955840 15936 10899636 13990 0 0 0 0
node "VSS" 81 122646 5268 10390 m2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 7756104 16428 794626 4030 112073122 106086 110747267 125354 15446591 30328 0 0 0 0
node "VDD" 214 94485.9 5485 7900 v2 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 7778407 24572 5663175 20848 88011407 88620 64944036 92864 31012240 26472 0 0 0 0
node "w_5404_4055#" 2160 110.16 5404 4055 nw 0 0 0 0 36720 772 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
substrate "VSUBS" 0 0 -1073741817 -1073741817 space 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
cap "VDD" "m1_5404_4055#" 2320.81
cap "VDD" "VN" 3797.94
cap "m2_2582_1554#" "VDD" 15.614
cap "VN" "VSS" 4767
cap "m2_1003_1555#" "m2_864_n933#" 43.3298
cap "m2_530_794#" "m2_864_n933#" 230.436
cap "m2_864_n933#" "VSS" 363.377
cap "m2_1498_1216#" "m2_864_n933#" 374.207
cap "VDD" "VO" 11351.1
cap "VO" "VSS" 15801.2
cap "m2_1003_1555#" "m2_530_794#" 368.324
cap "VDD" "m2_1003_1555#" 15.4514
cap "m2_1003_1555#" "VP" 78.232
cap "VDD" "IBIAS" 3797.94
cap "IBIAS" "VSS" 4767
cap "m1_5404_4055#" "VO" 4792.46
cap "m1_5404_4055#" "w_5404_4055#" 23.868
cap "m2_530_794#" "VP" 112.136
cap "VDD" "VSS" 31319
cap "VDD" "VP" 3797.94
cap "VP" "VSS" 4767
cap "m2_1498_1216#" "VSS" 363.377
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 51.3197
cap "CurrentMirror_layout_0/D3" "CurrentMirror_layout_0/S" 698.143
cap "CurrentMirror_layout_0/S" "CurrentMirror_layout_0/D1" 3.22744
cap "CurrentMirror_layout_0/D3" "CurrentMirror_layout_0/D1" 690.375
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" 262.005
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" 1610.1
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -246.231
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "VO" -527.1
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "VO" 2653.96
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "VO" -575.025
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "VO" 2653.96
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -101.02
cap "VO" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" -234.29
cap "CurrentMirror_layout_0/D1" "DiffPair_layout_0/w_n389_n527#" 284.196
cap "CurrentMirror_layout_0/D2" "CurrentMirror_layout_0/D1" 2100.43
cap "CurrentMirror_layout_0/D2" "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_3/a_50_n1050#" 2.27374e-13
cap "CurrentMirror_layout_0/D2" "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_0/a_n108_n1050#" 1.13687e-13
cap "CurrentMirror_layout_0/D2" "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_7/a_50_n1050#" 2.84217e-14
cap "CurrentMirror_layout_0/D2" "DiffPair_layout_0/w_n389_n527#" 704.237
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_9/a_50_n1050#" "CurrentMirror_layout_0/S" 87.2639
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_5/a_n50_n1076#" "CurrentMirror_layout_0/S" 3.22744
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_9/a_50_n1050#" "CurrentMirror_layout_0/D2" -2.84217e-14
cap "CurrentMirror_layout_0/sky130_fd_pr__nfet_01v8_RC9KLY_5/a_n50_n1076#" "CurrentMirror_layout_0/D2" -82.205
cap "VO" "CurrentMirror_layout_0/S" 77.5641
cap "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "m1_5404_4055#" 190.612
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/G1" 322.73
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 2.13163e-14
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/G1" 66.7336
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -98.6
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 1017.21
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_6/a_n50_n526#" 221.055
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_n50_n526#" 187.705
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_2/a_n50_n526#" 221.055
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/G1" -80.8235
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 401.3
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" 493.62
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 4.54747e-13
cap "DiffPair_layout_0/G1" "DiffPair_layout_0/D1" 51.65
cap "DiffPair_layout_0/w_n389_n527#" "m1_5404_4055#" 613.17
cap "PMOS2_0/S" "m1_5404_4055#" 38.8284
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 222.724
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_18/a_n50_n526#" 185.639
cap "m1_5404_4055#" "PMOS2_0/S" 5.3352
cap "PMOS2_0/S" "VO" 18.9696
cap "PMOS_Load_0/S" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 3.06
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -15.6202
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" -96.8202
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 7.8859
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" -315.819
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/w_n389_n527#" 322.73
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 90.195
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/G2" 214.483
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 216.993
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/G2" 89.92
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" -23.985
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_3/a_n50_n526#" 42.74
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/w_n389_n527#" 252.378
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" 36.485
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "PMOS_Load_0/S" 3.366
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/w_n389_n527#" 57.2455
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/G2" 111.527
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n50_n526#" -72.9359
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_7/a_n50_n526#" 42.74
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" 98.1339
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_0/a_n108_n500#" "PMOS_Load_0/S" 2.958
cap "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_1/a_50_n500#" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_3/a_n50_n526#" 52.3
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/D2" 252.378
cap "DiffPair_layout_0/D2" "PMOS_Load_0/S" 3.366
cap "DiffPair_layout_0/S" "DiffPair_layout_0/D2" 112.045
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/G2" -51
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/D2" -198.66
cap "DiffPair_layout_0/S" "DiffPair_layout_0/D1" -132.44
cap "DiffPair_layout_0/D2" "DiffPair_layout_0/G2" 216.912
cap "DiffPair_layout_0/w_n389_n527#" "m1_5404_4055#" 648.543
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/S" 472.795
cap "PMOS_Load_0/S" "DiffPair_layout_0/D1" 6.018
cap "PMOS_Load_0/S" "m1_5404_4055#" 58.641
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/D2" 223.993
cap "DiffPair_layout_0/D1" "DiffPair_layout_0/sky130_fd_pr__nfet_01v8_6YBK2C_19/a_n50_n526#" 16.85
cap "DiffPair_layout_0/w_n389_n527#" "DiffPair_layout_0/D1" 281.355
cap "DiffPair_layout_0/G2" "DiffPair_layout_0/D1" 315.028
cap "PMOS2_0/S" "m1_5404_4055#" 7.56
cap "PMOS2_0/D" "PMOS2_0/G" 897.876
cap "PMOS2_0/D" "PMOS2_0/S" 622.285
cap "PMOS2_0/S" "VO" -203.085
cap "PMOS_Load_0/D1" "PMOS_Load_0/S" -99.4994
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 786.318
cap "PMOS_Load_0/D2" "PMOS_Load_0/D1" 1139.21
cap "PMOS_Load_0/S" "PMOS_Load_0/D1" 126.929
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 200.884
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" "PMOS_Load_0/D2" 585.435
cap "PMOS_Load_0/D1" "PMOS_Load_0/D1" -73.68
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" 967.005
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" 172.201
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 384.612
cap "PMOS_Load_0/D1" "PMOS_Load_0/S" 337.38
cap "PMOS_Load_0/D1" "PMOS_Load_0/D2" -1.44
cap "PMOS2_0/S" "PMOS_Load_0/D2" 118.104
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n108_n600#" "PMOS_Load_0/S" 8.04255
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/S" 142.558
cap "PMOS_Load_0/D2" "PMOS_Load_0/S" 7.73381
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" 18.7864
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS_Load_0/S" 24.35
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/S" 1564.78
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_7/a_50_n600#" 8.80851
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_7/a_50_n600#" "PMOS_Load_0/D2" 5.68434e-14
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS_Load_0/S" 131.82
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" "PMOS_Load_0/S" 611.65
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_3/a_50_n600#" 8.80851
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n108_n600#" "PMOS_Load_0/D2" -82.205
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 413.144
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_0/a_n50_n626#" "PMOS_Load_0/D2" 268.73
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_3/a_50_n600#" "PMOS_Load_0/D2" -2.27374e-13
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" 39.2553
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_50_n600#" "PMOS_Load_0/D2" 155.002
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_12/a_n108_n600#" 8.80851
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/S" 1384.48
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_n50_n626#" 611.65
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_16/a_n108_n600#" "PMOS_Load_0/S" 8.80851
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_6/a_n50_n626#" "PMOS_Load_0/D2" 268.73
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 261.66
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS_Load_0/S" 49.32
cap "PMOS_Load_0/S" "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_19/a_50_n600#" 8.80851
cap "PMOS_Load_0/S" "PMOS_Load_0/D2" 56.54
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1384.48
cap "PMOS_Load_0/sky130_fd_pr__pfet_01v8_lvt_EEU9S7_15/a_n50_n626#" "PMOS_Load_0/S" 215.825
cap "PMOS_Load_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -12.32
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS2_0/S" -206.885
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS2_0/S" -14.85
cap "PMOS2_0/S" "PMOS_Load_0/D2" 175.002
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 57.5463
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "PMOS2_0/S" 1261.4
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 49.32
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1384.48
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1384.48
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 49.32
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1204.02
cap "PMOS2_0/S" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" 63.55
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "PMOS2_0/S" -1352.34
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 117.549
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 386.26
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 154
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 4067.93
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "VDD" -1378.37
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "VDD" -1262.8
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "VDD" -870.93
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 253.499
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "VDD" 1486.5
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 263.284
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 253.499
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 2470.58
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "VDD" -1262.8
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" -1262.8
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 3985.43
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "VDD" -1240.4
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 4239.25
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 453.67
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 70.11
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 518.775
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 1645.15
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" 386.8
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 2187.5
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 2443
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 2538.14
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 92.9015
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" 854.147
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 1561.69
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 2443
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 2443
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" 2241.96
cap "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "VDD" 1111.78
cap "VDD" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" -70.3871
merge "PMOS_Load_0/D1" "DiffPair_layout_0/D1" -1862.94 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -138970 -1328 -373736 -3878 0 0 0 0 0 0
merge "DiffPair_layout_0/D1" "m2_3531_794#"
merge "m2_3531_794#" "m2_530_794#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/m3_n3150_n1100#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/VSUBS" -11197.3 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -5394990 -20718 0 0 0 0 0 0 -777170 -11492 0 0 0 0
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/VSUBS" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/VSUBS"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/VSUBS" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/m3_n3150_n1100#" "PMOS_Load_0/VSUBS"
merge "PMOS_Load_0/VSUBS" "PMOS2_0/VSUBS"
merge "PMOS2_0/VSUBS" "DiffPair_layout_0/w_n389_n527#"
merge "DiffPair_layout_0/w_n389_n527#" "CurrentMirror_layout_0/S"
merge "CurrentMirror_layout_0/S" "VSS"
merge "VSS" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/VSUBS"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/VSUBS" "VSUBS"
merge "PMOS2_0/G" "PMOS_Load_0/D2" -4296.62 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 3335 -472 -935032 -2260 48840 -2230 0 0 0 0 0 0
merge "PMOS_Load_0/D2" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/c1_n2450_n2400#" "m1_5404_4055#"
merge "m1_5404_4055#" "DiffPair_layout_0/D2"
merge "DiffPair_layout_0/D2" "m2_2582_1554#"
merge "m2_2582_1554#" "m2_1003_1555#"
merge "DiffPair_layout_0/S" "CurrentMirror_layout_0/D2" -2812.1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -24247 -2740 -306139 -6596 0 0 0 0 0 0
merge "CurrentMirror_layout_0/D2" "m2_1498_1216#"
merge "m2_1498_1216#" "m2_864_n933#"
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_1/c1_n3050_n1000#" "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" -38606 0 0 0 0 -26690 -772 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -605657 -26722 1466048 -14587 -26748840 -32187 -2287682 -27214 -21157388 -26923 0 0 0 0
merge "sky130_fd_pr__cap_mim_m3_1_N3PKNJ_0/c1_n3050_n1000#" "PMOS2_0/S"
merge "PMOS2_0/S" "w_5404_4055#"
merge "w_5404_4055#" "PMOS_Load_0/S"
merge "PMOS_Load_0/S" "VDD"
merge "PMOS2_0/D" "CurrentMirror_layout_0/D3" -11123.1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -4857782 -20481 -3468453 -7600 -654505 -20469 0 0 0 0
merge "CurrentMirror_layout_0/D3" "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#"
merge "sky130_fd_pr__cap_mim_m3_1_TQVBRR_0/m3_n2550_n2500#" "VO"
merge "DiffPair_layout_0/G1" "VN" 170.229 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 161075 -328 167475 0 0 0 0 0 0 0 0 0
merge "DiffPair_layout_0/G2" "VP" -475.348 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -26880 -1166 0 0 0 0 0 0 0 0 0 0
merge "CurrentMirror_layout_0/D1" "IBIAS" -476.836 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 -452007 -342 0 0 0 0 0 0 0 0
                                                                                                                                                n0 VSS VSS nch w=0.39u l=0.06u
MU1_7-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_0-M_u4 n0 A1 VSS VSS nch w=0.195u l=0.06u
M_u7_0-M_u3 n0 A2 VSS VSS nch w=0.195u l=0.06u
M_u7_1-M_u4 n0 A1 VSS VSS nch w=0.195u l=0.06u
M_u7_1-M_u3 n0 A2 VSS VSS nch w=0.195u l=0.06u
M_u7_2-M_u4 n0 A1 VSS VSS nch w=0.195u l=0.06u
M_u7_2-M_u3 n0 A2 VSS VSS nch w=0.195u l=0.06u
MU1_0-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_1-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_2-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_3-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_4-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_5-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_6-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
MU1_7-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_0-M_u1 X_u7_0-net8 A2 VDD VDD pch w=0.52u l=0.06u
M_u7_0-M_u2 n0 A1 X_u7_0-net8 VDD pch w=0.52u l=0.06u
M_u7_1-M_u1 X_u7_1-net8 A2 VDD VDD pch w=0.52u l=0.06u
M_u7_1-M_u2 n0 A1 X_u7_1-net8 VDD pch w=0.52u l=0.06u
M_u7_2-M_u1 X_u7_2-net8 A2 VDD VDD pch w=0.52u l=0.06u
M_u7_2-M_u2 n0 A1 X_u7_2-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt OR2XD1 A1 A2 Z VDD VSS
MU1-M_u2 Z net7 VSS VSS nch w=0.39u l=0.06u
M_u7-M_u4 net7 A1 VSS VSS nch w=0.39u l=0.06u
M_u7-M_u3 net7 A2 VSS VSS nch w=0.39u l=0.06u
MU1-M_u3 Z net7 VDD VDD pch w=0.52u l=0.06u
M_u7-M_u1 X_u7-net8 A2 VDD VDD pch w=0.52u l=0.06u
M_u7-M_u2 net7 A1 X_u7-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt OR3D0 A1 A2 A3 Z VDD VSS
M_u4-M_u2 Z net7 VSS VSS nch w=0.195u l=0.06u
MU42-M_u6 net7 A3 VSS VSS nch w=0.195u l=0.06u
MU42-M_u5 net7 A2 VSS VSS nch w=0.195u l=0.06u
MU42-M_u4 net7 A1 VSS VSS nch w=0.195u l=0.06u
M_u4-M_u3 Z net7 VDD VDD pch w=0.26u l=0.06u
MU42-M_u1 XU42-net9 A1 VDD VDD pch w=0.26u l=0.06u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD pch w=0.26u l=0.06u
MU42-M_u3 net7 A3 XU42-net12 VDD pch w=0.26u l=0.06u
.ends
.subckt OR3D1 A1 A2 A3 Z VDD VSS
M_u4-M_u2 Z net7 VSS VSS nch w=0.39u l=0.06u
MU42-M_u6 net7 A3 VSS VSS nch w=0.195u l=0.06u
MU42-M_u5 net7 A2 VSS VSS nch w=0.195u l=0.06u
MU42-M_u4 net7 A1 VSS VSS nch w=0.195u l=0.06u
M_u4-M_u3 Z net7 VDD VDD pch w=0.52u l=0.06u
MU42-M_u1 XU42-net9 A1 VDD VDD pch w=0.52u l=0.06u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD pch w=0.52u l=0.06u
MU42-M_u3 net7 A3 XU42-net12 VDD pch w=0.52u l=0.06u
.ends
.subckt OR3D2 A1 A2 A3 Z VDD VSS
M_u4_0-M_u2 Z net12 VSS VSS nch w=0.39u l=0.06u
M_u4_1-M_u2 Z net12 VSS VSS nch w=0.39u l=0.06u
MU42-M_u6 net12 A3 VSS VSS nch w=0.195u l=0.06u
MU42-M_u5 net12 A2 VSS VSS nch w=0.195u l=0.06u
MU42-M_u4 net12 A1 VSS VSS nch w=0.195u l=0.06u
M_u4_0-M_u3 Z net12 VDD VDD pch w=0.52u l=0.06u
M_u4_1-M_u3 Z net12 VDD VDD pch w=0.52u l=0.06u
MU42-M_u1 XU42-net9 A1 VDD VDD pch w=0.52u l=0.06u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD pch w=0.52u l=0.06u
MU42-M_u3 net12 A3 XU42-net12 VDD pch w=0.52u l=0.06u
.ends
.subckt OR3D4 A1 A2 A3 Z VDD VSS
M_u4_0-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_1-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_2-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_3-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU42_0-M_u6 p0 A3 VSS VSS nch w=0.195u l=0.06u
MU42_0-M_u5 p0 A2 VSS VSS nch w=0.195u l=0.06u* NGSPICE file created from OpampM_PL.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_RC9KLY a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS
X0 a_50_n1050# a_n50_n1076# a_n108_n1050# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=500000u
.ends

.subckt CurrentMirror_layout D3 D2 D1 S
Xsky130_fd_pr__nfet_01v8_RC9KLY_1 D2 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_3 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_2 S D1 D2 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_4 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_5 D1 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_6 S D1 D1 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_7 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_8 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_9 D3 D1 S S sky130_fd_pr__nfet_01v8_RC9KLY
Xsky130_fd_pr__nfet_01v8_RC9KLY_0 S D1 D3 S sky130_fd_pr__nfet_01v8_RC9KLY
.ends

.subckt sky130_fd_pr__nfet_01v8_6YBK2C a_50_n500# a_n50_n526# a_n108_n500# VSUBS
X0 a_50_n500# a_n50_n526# a_n108_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt DiffPair_layout D2 D1 G2 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
Xsky130_fd_pr__nfet_01v8_6YBK2C_10 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_11 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_13 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_12 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_14 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_15 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_16 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_17 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_18 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_19 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_0 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_2 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_1 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_3 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_4 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_5 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_6 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_7 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_8 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_9 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_EEU9S7 w_n144_n662# a_50_n600# a_n50_n626#
+ a_n108_n600# VSUBS
X0 a_50_n600# a_n50_n626# a_n108_n600# w_n144_n662# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
.ends

.subckt PMOS_Load D2 D1 S VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_0 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_1 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_10 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_2 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_11 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_3 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_12 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_4 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_13 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_5 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_14 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_7 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_6 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_15 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_8 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_16 S S D1 D1 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_9 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_17 S D2 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_19 S D1 D1 S VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
Xsky130_fd_pr__pfet_01v8_lvt_EEU9S7_18 S S D1 D2 VSUBS sky130_fd_pr__pfet_01v8_lvt_EEU9S7
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TQVBRR m3_n2550_n2500# c1_n2450_n2400# VSUBS
X0 c1_n2450_n2400# m3_n2550_n2500# sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.4e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_N3PKNJ c1_n3050_n1000# m3_n3150_n1100# VSUBS
X0 c1_n3050_n1000# m3_n3150_n1100# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_WFBLZ7 a_50_n1420# a_n50_n1446# w_n144_n1482# a_n108_n1420#
+ VSUBS
X0 a_50_n1420# a_n50_n1446# a_n108_n1420# w_n144_n1482# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.42e+07u l=500000u
.ends

.subckt PMOS2 G D S VSUBS
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_19 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_0 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_1 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_2 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_3 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_5 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_4 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_6 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_7 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_8 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_9 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_20 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_21 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_10 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_22 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_11 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_23 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_12 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_24 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_13 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_14 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_15 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_16 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_17 S G S D VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
Xsky130_fd_pr__pfet_01v8_lvt_WFBLZ7_18 D G S S VSUBS sky130_fd_pr__pfet_01v8_lvt_WFBLZ7
.ends

.subckt OpampM_PL VSS VDD VO VP VN IBIAS
XCurrentMirror_layout_0 VO DiffPair_layout_0/S IBIAS VSS CurrentMirror_layout
XDiffPair_layout_0 PMOS2_0/G PMOS_Load_0/D1 VP VN DiffPair_layout_0/S VSS DiffPair_layout
XPMOS_Load_0 PMOS2_0/G PMOS_Load_0/D1 VDD VSS PMOS_Load
Xsky130_fd_pr__cap_mim_m3_1_TQVBRR_0 VO PMOS2_0/G VSS sky130_fd_pr__cap_mim_m3_1_TQVBRR
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_0 VDD VSS VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
Xsky130_fd_pr__cap_mim_m3_1_N3PKNJ_1 VDD VSS VSS sky130_fd_pr__cap_mim_m3_1_N3PKNJ
XPMOS2_0 PMOS2_0/G VO VDD VSS PMOS2
.ends

                                                                                                                                                                         l=0.06u
MI165 net63 CDN VSS VSS nch w=0.15u l=0.06u
MI164 net82 d1 net63 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net82 VSS nch w=0.15u l=0.06u
MI169 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI161 net67 SI VSS VSS nch w=0.15u l=0.06u
MI160 net177 SE net67 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.39u l=0.06u
MI166-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI151-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q net0140 VSS VSS nch w=0.39u l=0.06u
MI174-M_u2 net62 net0140 VSS VSS nch w=0.23u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI32-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI158-M_u4 XI158-net6 CDN VSS VSS nch w=0.35u l=0.06u
MI158-M_u3 net0140 net163 XI158-net6 VSS nch w=0.35u l=0.06u
MI166-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI151-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 Q net0140 VDD VDD pch w=0.52u l=0.06u
MI174-M_u3 net62 net0140 VDD VDD pch w=0.52u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI32-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI155 net62 INCP net163 VDD pch w=0.16u l=0.06u
MI170 net132 SE net69 VDD pch w=0.44u l=0.06u
MI163 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI162 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net132 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net132 VDD pch w=0.29u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 INCPB net163 VDD pch w=0.29u l=0.06u
MI158-M_u2 net0140 CDN VDD VDD pch w=0.44u l=0.06u
MI158-M_u1 net0140 net163 VDD VDD pch w=0.44u l=0.06u
.ends
.subckt SDFCND2 SI D SE CP CDN Q QN VDD VSS
MI150 net62 INCPB d2 VSS nch w=0.15u l=0.06u
MI149 d1 INCP d2 VSS nch w=0.2u l=0.06u
MI165 net63 CDN VSS VSS nch w=0.15u l=0.06u
MI164 net82 d1 net63 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net82 VSS nch w=0.15u l=0.06u
MI169 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI161 net67 SI VSS VSS nch w=0.15u l=0.06u
MI160 net177 SE net67 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.39u l=0.06u
MI178-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI179-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI171-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI172-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI151-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI176-M_u2 net62 d3 VSS VSS nch w=0.21u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI158_0-M_u4 XI158_0-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_0-M_u3 d3 d2 XI158_0-net6 VSS nch w=0.23u l=0.06u
MI158_1-M_u4 XI158_1-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_1-M_u3 d3 d2 XI158_1-net6 VSS nch w=0.23u l=0.06u
MI178-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI179-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI171-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI172-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI151-M_u3 QN net62 VDputs stdout "Sourcing design .magicrc for technology sky130A ..."

# Put grid on 0.005 pitch.  This is important, as some commands don't
# rescale the grid automatically (such as lef read?).

set scalefac [tech lambda]
if {[lindex $scalefac 1] < 2} {
    scalegrid 1 2
}

# drc off
drc euclidean on
# Change this to a fixed number for repeatable behavior with GDS writes
# e.g., "random seed 12345"
catch {random seed}

# Turn off the scale option on ext2spice or else it conflicts with the
# scale in the model files.
ext2spice scale off

# Allow override of PDK path from environment variable PDKPATH
if {[catch {set PDKPATH $env(PDKPATH)}]} {
    set PDKPATH "/home/shahid/SkywaterPDK//sky130A"
}

# loading technology
tech load $PDKPATH/libs.tech/magic/sky130A.tech

# load device generator
source $PDKPATH/libs.tech/magic/sky130A.tcl

# load bind keys (optional)
# source $PDKPATH/libs.tech/magic/sky130A-BindKeys

# set units to lambda grid 
snap lambda

# set sky130 standard power, ground, and substrate names
set VDD VPWR
set GND VGND
set SUB VSUBS

# Allow override of type of magic library views used, "mag" or "maglef",
# from environment variable MAGTYPE

if {[catch {set MAGTYPE $env(MAGTYPE)}]} {
   set MAGTYPE mag
}

# add path to reference cells
if {[file isdir ${PDKPATH}/libs.ref/${MAGTYPE}]} {
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_pr
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_io
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_hd
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_hdll
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_hs
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_hvl
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_lp
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_ls
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_fd_sc_ms
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_osu_sc
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_osu_sc_t18
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_ml_xx_hd
    addpath ${PDKPATH}/libs.ref/${MAGTYPE}/sky130_sram_macros
} else {
    addpath ${PDKPATH}/libs.ref/sky130_fd_pr/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_io/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_hd/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_hdll/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_hs/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_hvl/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_lp/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_ls/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_fd_sc_ms/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_osu_sc/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_osu_sc_t18/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_ml_xx_hd/${MAGTYPE}
    addpath ${PDKPATH}/libs.ref/sky130_sram_macros/${MAGTYPE}
}

# add path to GDS cells

# add path to IP from catalog.  This procedure defined in the PDK script.
catch {magic::query_mylib_ip}
# add path to local IP from user design space.  Defined in the PDK script.
catch {magic::query_my_projects}
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      111 SE VSS VSS nch w=0.15u l=0.06u
MI32-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI26 net161 d3 VSS VSS nch w=0.15u l=0.06u
MI149 d1 INCP d2 VSS nch w=0.2u l=0.06u
MI29 d2 INCPB net161 VSS nch w=0.15u l=0.06u
MI165 net63 CDN VSS VSS nch w=0.15u l=0.06u
MI164 net82 d1 net63 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net82 VSS nch w=0.15u l=0.06u
MI169 net177 D net0103 VSS nch w=0.26u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI161 net67 SI VSS VSS nch w=0.15u l=0.06u
MI160 net177 SE net67 VSS nch w=0* NGSPICE file created from DiffPair_layout.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_6YBK2C a_50_n500# a_n50_n526# a_n108_n500# VSUBS
X0 a_50_n500# a_n50_n526# a_n108_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends


* Top level circuit DiffPair_layout

Xsky130_fd_pr__nfet_01v8_6YBK2C_10 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_11 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_13 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_12 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_14 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_15 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_16 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_17 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_18 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_19 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS
+ sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_0 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_2 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_1 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_3 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_4 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_5 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_6 S G2 D2 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_7 D1 G1 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_8 S G1 D1 sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
Xsky130_fd_pr__nfet_01v8_6YBK2C_9 D2 G2 S sky130_fd_pr__nfet_01v8_6YBK2C_9/VSUBS sky130_fd_pr__nfet_01v8_6YBK2C
.end

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       et177 SE net67 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.39u l=0.06u
MI29 d2 INCPB net078 VSS nch w=0.15u l=0.06u
MI178-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI171-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI172-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI158_0-M_u4 XI158_0-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_0-M_u3 d3 d2 XI158_0-net6 VSS nch w=0.23u l=0.06u
MI158_1-M_u4 XI158_1-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_1-M_u3 d3 d2 XI158_1-net6 VSS nch w=0.23u l=0.06u
MI178-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI171-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI172-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI152-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI28 d2 INCP net0119 VDD pch w=0.15u l=0.06u
MI24 net0119 d3 VDD VDD pch w=0.15u l=0.06u
MI170 net132 SE net69 VDD pch w=0.44u l=0.06u
MI175 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI162 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net132 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net132 VDD pch w=0.29u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI174 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 INCPB d2 VDD pch w=0.29u l=0.06u
MI158_0-M_u2 d3 CDN VDD VDD pch w=0.52u l=0.06u
MI158_0-M_u1 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI158_1-M_u2 d3 CDN VDD VDD pch w=0.52u l=0.06u
MI158_1-M_u1 d3 d2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFCNQD4 SI D SE CP CDN Q VDD VSS
MI149 d1 INCP d2 VSS nch w=0.2u l=0.06u
MI26 net090 d3 VSS VSS nch w=0.15u l=0.06u
MI165 net63 CDN VSS VSS nch w=0.15u l=0.06u
MI164 net82 d1 net63 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net82 VSS nch w=0.15u l=0.06u
MI169 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI77 d0 net0112 net177 VSS nch w=0.3u l=0.06u
MI161 net67 SI VSS VSS nch w=0.15u l=0.06u
MI160 net177 SE net67 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.39u l=0.06u
MI29 d2 net0112 net090 VSS nch w=0.15u l=0.06u
MI167-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI185-M_u2 net0112 CP VSS VSS nch w=0.39u l=0.06u
MI186-M_u2 INCP net0112 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI176-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI177-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI158_0-M_u4 XI158_0-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_0-M_u3 d3 d2 XI158_0-net6 VSS nch w=0.23u l=0.06u
MI158_1-M_u4 XI158_1-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158_1-M_u3 d3 d2 XI158_1-net6 VSS nch w=0.23u l=0.06u
MI167-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI185-M_u3 net0112 CP VDD VDD pch w=0.52u l=0.06u
MI186-M_u3 INCP net0112 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI176-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI177-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI28 d2 INCP net0135 VDD pch w=0.15u l=0.06u
MI24 net0135 d3 VDD VDD pch w=0.15u l=0.06u
MI170 net132 SE net69 VDD pch w=0.44u l=0.06u
MI175 d0 net0112 net166 VDD pch w=0.15u l=0.06u
MI162 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net132 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net132 VDD pch w=0.29u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI174 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 net0112 d2 VDD pch w=0.29u l=0.06u
MI158_0-M_u2 d3 CDN VDD VDD pch w=0.52u l=0.06u
MI158_0-M_u1 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI158_1-M_u2 d3 CDN VDD VDD pch w=0.52u l=0.06u
MI158_1-M_u1 d3 d2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFCSND0 SI D SE CP CDN SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 D net0102 VSS nch w=0.26u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net0102 net0108 VSS VSS nch w=0.26u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net0108 SE VSS VSS nch w=0.15u l=0.06u
MI104-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net0108 SE VDD VDD pch w=0.2u l=0.06u
MI104-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI102 net104 D net107 VDD pch w=0.33u l=0.06u
MI45 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net0108 net148 VDD pch w=0.15u l=0.06u
MI73 net107 SE VDD VDD pch w=0.33u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net148 SI VDD VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSND1 SI D SE CP CDN SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.35u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI32-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI32-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI102 net104 SE net107 VDD pch w=0.44u l=0.06u
MI104 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSND2 SI D SE CP CDN SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.35u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI100-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI106-M_u4 XI106-net6 d3 VSS VSS nch w=0.35u l=0.06u
MI106-M_u3 d4 SDN XI106-net6 VSS nch w=0.35u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI100-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI108-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI102 net104 SE net107 VDD pch w=0.44u l=0.06u
MI45 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI106-M_u2 d4 d3 VDD VDD pch w=0.38u l=0.06u
MI106-M_u1 d4 SDN VDD VDD pch w=0.38u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSND4 SI D SE CP CDN SDN Q QN VDD VSS
MI91 d4 net0120 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.35u l=0.06u
MI77 d0 net0120 net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI114-M_u2 INCP net0120 VSS VSS nch w=0.39u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI100-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI107-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI109-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI110-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI113-M_u2 net0120 CP VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI106-M_u4 XI106-net6 d3 VSS VSS nch w=0.35u l=0.06u
MI106-M_u3 d4 SDN XI106-net6 VSS nch w=0.35u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.17u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.17u l=0.06u
MI105-M_u4 XI105-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI105-M_u3 d3 CDN XI105-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI114-M_u3 INCP net0120 VDD VDD pch w=0.52u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI100-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI107-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI108-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI109-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI110-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI113-M_u3 net0120 CP VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI102 net104 SE net107 VDD pch w=0.44u l=0.06u
MI45 d0 net0120 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 net0120 d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI106-M_u2 d4 d3 VDD VDD pch w=0.38u l=0.06u
MI106-M_u1 d4 SDN VDD VDD pch w=0.38u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI105-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI105-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSNQD0 SI D SE CP CDN SDN Q VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 D net0102 VSS nch w=0.26u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net0102 net0108 VSS VSS nch w=0.26u l=0.06u
MI105-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net0108 SE VSS VSS nch w=0.15u l=0.06u
MI31-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.34u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.34u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI105-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net0108 SE VDD VDD pch w=0.2u l=0.06u
MI31-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI102 net104 D net107 VDD pch w=0.33u l=0.06u
MI45 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net0108 net148 VDD pch w=0.15u l=0.06u
MI73 net107 SE VDD VDD pch w=0.33u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net148 SI VDD VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSNQD1 SI D SE CP CDN SDN Q VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.39u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI31-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI103-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.2u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.2u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI31-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI103-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI102 net104 SE net107 VDD pch w=0.4u l=0.06u
MI105 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.49u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.32u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.2u l=0.06u
MI104 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.15u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.15u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSNQD2 SI D SE CP CDN SDN Q VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.39u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI107-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI106-M_u4 XI106-net6 d2 VSS VSS nch w=0.17u l=0.06u
MI106-M_u3 d3 CDN XI106-net6 VSS nch w=0.17u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.15u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.15u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI107-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI102 net104 SE net107 VDD pch w=0.4u l=0.06u
MI45 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.49u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.32u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI106-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI106-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.15u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.15u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFCSNQD4 SI D SE CP CDN SDN Q VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCP net86 VSS nch w=0.15u l=0.06u
MI101 net177 net120 net107 VSS nch w=0.39u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.3u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net107 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI104-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI32-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.15u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.15u l=0.06u
MI106-M_u4 XI106-net6 d2 VSS VSS nch w=0.19u l=0.06u
MI106-M_u3 d3 CDN XI106-net6 VSS nch w=0.19u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.32u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.32u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI108-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI104-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI32-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI102 net104 SE net107 VDD pch w=0.4u l=0.06u
MI45 d0 INCPB net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net107 D VDD VDD pch w=0.49u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.32u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.15u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.15u l=0.06u
MI106-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI106-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFD0 SI D SE CP Q QN VDD VSS
MI39 net37 D net64 VSS nch w=0.26u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 INCPB d2 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.16u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 net57 VSS VSS nch w=0.26u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.195u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI41-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.26u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI41-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCP d2 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net0111 SE VDD VDD pch w=0.33u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 D net0111 VDD pch w=0.33u l=0.06u
.ends
.subckt SDFD1 SI D SE CP Q QN VDD VSS
MI39 net37 net57 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 INCPB d2 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.18u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.195u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI41-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=0.26u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI41-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCP d2 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFD2 SI D SE CP Q QN VDD VSS
MI39 net37 net57 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 INCPB d2 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.16u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI38-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI43-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI38-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI43-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCP d2 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFD4 SI D SE CP Q QN VDD VSS
MI39 net37 net0139 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 INCPB d2 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.19u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI38-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.78u l=0.06u
MI44-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI45-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI46-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI47-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI49-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI50-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net0139 SE VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI38-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=1.04u l=0.06u
MI44-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI45-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI46-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI47-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI49-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI50-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net0139 SE VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCP d2 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net0139 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFKCND0 SI D SE CP CN Q QN VDD VSS
MI138-M_u2 QN net69 VSS VSS nch w=0.195u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI139-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.15u l=0.06u
MI140-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI142-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.195u l=0.06u
MI80 net135 D VSS VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 QN net69 VDD VDD pch w=0.26u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI139-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.2u l=0.06u
MI140-M_u3 net93 net155 VDD VDD pch w=0.295u l=0.06u
MI142-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.2u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.495u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.26u l=0.06u
MI77 VDD D net132 VDD pch w=0.26u l=0.06u
.ends
.subckt SDFKCND1 SI D SE CP CN Q QN VDD VSS
MI138-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI144-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI143-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI141-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.33u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.39u l=0.06u
MI80 net135 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI144-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI143-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI141-M_u3 net93 net155 VDD VDD pch w=0.295u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.495u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCND2 SI D SE CP CN Q QN VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI142-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 p0 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.33u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB p0 VSS nch w=0.27u l=0.06u
MI101 p0 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.39u l=0.06u
MI80 net135 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI142-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 p0 VDD VDD pch w=0.295u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.495u l=0.06u
MI127 net109 INCP p0 VDD pch w=0.34u l=0.06u
MI99 p0 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCND4 SI D SE CP CN Q QN VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI145-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI49-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI42_0-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI42_1-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI141-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI146-M_u2 net69 net105 VSS VSS nch w=0.235u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI142-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI143-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI144-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.565u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.33u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.39u l=0.06u
MI80 net135 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI145-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI49-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI42_0-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI42_1-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI141-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI146-M_u3 net69 net105 VDD VDD pch w=0.315u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI142-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI143-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI144-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCNQD0 SI D SE CP CN Q VDD VSS
MI112 net93 INCP net71 VSS nch w=0.18u l=0.06u
MI122 net068 Q VSS VSS nch w=0.15u l=0.06u
MI64 net76 net85 VSS VSS nch w=0.195u l=0.06u
MI65 net146 net81 net76 VSS nch w=0.195u l=0.06u
MI62 net146 SE net101 VSS nch w=0.15u l=0.06u
MI121 net71 INCPB net068 VSS nch w=0.15u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI83 net155 INCPB net146 VSS nch w=0.23u l=0.06u
MI63 net101 net0106 VSS VSS nch w=0.15u l=0.06u
MI79 net81 CN net135 VSS nch w=0.15u l=0.06u
MI80 net135 D VSS VSS nch w=0.15u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net85 SE VSS VSS nch w=0.195u l=0.06u
MI126-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI127-M_u2 net0106 SI VSS VSS nch w=0.15u l=0.06u
MI129-M_u2 Q net71 VSS VSS nch w=0.39u l=0.06u
MI128-M_u2 net93 net155 VSS VSS nch w=0.34u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI45-M_u3 net85 SE VDD VDD pch w=0.29u l=0.06u
MI126-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI127-M_u3 net0106 SI VDD VDD pch w=0.15u l=0.06u
MI129-M_u3 Q net71 VDD VDD pch w=0.52u l=0.06u
MI128-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI50 net127 SE VDD VDD pch w=0.235u l=0.06u
MI82 net155 INCP net117 VDD pch w=0.3u l=0.06u
MI123 net71 INCP net0116 VDD pch w=0.15u l=0.06u
MI53 net117 net85 net139 VDD pch w=0.15u l=0.06u
MI51 net117 net81 net127 VDD pch w=0.235u l=0.06u
MI52 net139 net0106 VDD VDD pch w=0.15u l=0.06u
MI124 net0116 Q VDD VDD pch w=0.15u l=0.06u
MI119 net93 INCPB net71 VDD pch w=0.43u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI74 VDD CN net81 VDD pch w=0.2u l=0.06u
MI77 VDD D net81 VDD pch w=0.2u l=0.06u
.ends
.subckt SDFKCNQD1 SI D SE CP CN Q VDD VSS
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI139-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI140-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.33u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.39u l=0.06u
MI80 net135 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI139-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.295u l=0.06u
MI140-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.495u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCNQD2 SI D SE CP CN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI140-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.33u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.39u l=0.06u
MI80 net135 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.295u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.495u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCNQD4 SI D SE CP CN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.24u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI42_0-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI42_1-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI142-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.565u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.35u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 CN net135 VSS nch w=0.41u l=0.06u
MI80 net135 D VSS VSS nch w=0.41u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.52u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI42_0-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI42_1-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI142-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.51u l=0.06u
MI77 VDD D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKCSND0 SI D SE CP CN SN Q QN VDD VSS
MI140-M_u2 QN net69 VSS VSS nch w=0.195u l=0.06u
MI142-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.15u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI143-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI72-M_u2 net120 SN VSS VSS nch w=0.15u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI80 net91 CN VSS VSS nch w=0.195u l=0.06u
MI78 net132 net120 net91 VSS nch w=0.195u l=0.06u
MI79 net132 D net91 VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.26u l=0.06u
MI142-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.2u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.305u l=0.06u
MI143-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI72-M_u3 net120 SN VDD VDD pch w=0.2u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI77 net143 D net132 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.485u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.26u l=0.06u
MI75 VDD net120 net143 VDD pch w=0.27u l=0.06u
.ends
.subckt SDFKCSND1 SI D SE CP CN SN Q QN VDD VSS
MI138-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net120 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI80 net91 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net120 net91 VSS nch w=0.2u l=0.06u
MI79 net132 D net91 VSS nch w=0.2u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.305u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net120 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI77 net143 D net132 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.485u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
MI75 VDD net120 net143 VDD pch w=0.27u l=0.06u
.ends
.subckt SDFKCSND2 SI D SE CP CN SN Q QN VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI142-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI141-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI139-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net127 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D net104 VSS nch w=0.2u l=0.06u
MI80 net104 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net127 net104 VSS nch w=0.2u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI142-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI141-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.305u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net127 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI75 VDD net127 net151 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.485u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI77 net151 D net132 VDD pch w=0.27u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
.ends
.subckt SDFKCSND4 SI D SE CP CN SN Q QN VDD VSS
MI142-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI147-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI141-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI139-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.42u l=0.06u
MI143-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.235u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI144-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI145-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI146-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net127 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.565u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D net104 VSS nch w=0.2u l=0.06u
MI80 net104 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net127 net104 VSS nch w=0.2u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI142-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI147-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI141-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.68u l=0.06u
MI143-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.315u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI144-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI145-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI146-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net127 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI75 VDD net127 net151 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI77 net151 D net132 VDD pch w=0.27u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
.ends
.subckt SDFKCSNQD0 SI D SE CP CN SN Q VDD VSS
MI131 net80 net85 VSS VSS nch w=0.175u l=0.06u
MI130 net146 net81 net80 VSS nch w=0.175u l=0.06u
MI132 net146 SE net65 VSS nch w=0.15u l=0.06u
MI118 net93 INCP net74 VSS nch w=0.21u l=0.06u
MI95 net161 INCP net104 VSS nch w=0.15u l=0.06u
MI135 net74 INCPB net074 VSS nch w=0.15u l=0.06u
MI122 net074 Q VSS VSS nch w=0.15u l=0.06u
MI83 net161 INCPB net146 VSS nch w=0.23u l=0.06u
MI133 net65 net0110 VSS VSS nch w=0.15u l=0.06u
MI96 net104 net93 VSS VSS nch w=0.15u l=0.06u
MI78 net81 net83 net135 VSS nch w=0.195u l=0.06u
MI79 net81 D net135 VSS nch w=0.195u l=0.06u
MI80 net135 CN VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net85 SE VSS VSS nch w=0.195u l=0.06u
MI141-M_u2 net0110 SI VSS VSS nch w=0.15u l=0.06u
MI121-M_u2 Q net74 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 net161 VSS VSS nch w=0.34u l=0.06u
MI140-M_u2 net83 SN VSS VSS nch w=0.15u l=0.06u
MI139-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI45-M_u3 net85 SE VDD VDD pch w=0.26u l=0.06u
MI141-M_u3 net0110 SI VDD VDD pch w=0.15u l=0.06u
MI121-M_u3 Q net74 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 net161 VDD VDD pch w=0.34u l=0.06u
MI140-M_u3 net83 SN VDD VDD pch w=0.2u l=0.06u
MI126 net117 net81 net140 VDD pch w=0.255u l=0.06u
MI82 net161 INCP net117 VDD pch w=0.3u l=0.06u
MI128 net117 net85 net129 VDD pch w=0.2u l=0.06u
MI127 net140 SE VDD VDD pch w=0.255u l=0.06u
MI129 net129 net0110 VDD VDD pch w=0.2u l=0.06u
MI136 net0126 Q VDD VDD pch w=0.15u l=0.06u
MI123 net74 INCP net0126 VDD pch w=0.15u l=0.06u
MI125 net93 INCPB net74 VDD pch w=0.43u l=0.06u
MI74 VDD CN net81 VDD pch w=0.375u l=0.06u
MI94 net170 net93 VDD VDD pch w=0.15u l=0.06u
MI93 net161 INCPB net170 VDD pch w=0.15u l=0.06u
MI75 VDD net83 net173 VDD pch w=0.375u l=0.06u
MI77 net173 D net81 VDD pch w=0.375u l=0.06u
.ends
.subckt SDFKCSNQD1 SI D SE CP CN SN Q VDD VSS
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI139-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI140-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net120 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI80 net91 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net120 net91 VSS nch w=0.2u l=0.06u
MI79 net132 D net91 VSS nch w=0.2u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI139-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI140-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.305u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net120 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI77 net143 D net132 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.485u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
MI75 VDD net120 net143 VDD pch w=0.27u l=0.06u
.ends
.subckt SDFKCSNQD2 SI D SE CP CN SN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI142-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI141-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI143-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net127 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.235u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D net104 VSS nch w=0.2u l=0.06u
MI80 net104 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net127 net104 VSS nch w=0.2u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI142-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI141-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.305u l=0.06u
MI143-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net127 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI75 VDD net127 net151 VDD pch w=0.27u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.485u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI77 net151 D net132 VDD pch w=0.27u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
.ends
.subckt SDFKCSNQD4 SI D SE CP CN SN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI146-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.365u l=0.06u
MI49-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.185u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI42_0-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI42_1-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net239 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.565u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI80 net216 CN VSS VSS nch w=0.2u l=0.06u
MI78 net132 net239 net216 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI79 net132 D net216 VSS nch w=0.2u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI146-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.515u l=0.06u
MI49-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI42_0-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI42_1-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net239 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.28u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI77 net271 D net132 VDD pch w=0.27u l=0.06u
MI74 VDD CN net132 VDD pch w=0.235u l=0.06u
MI75 VDD net239 net271 VDD pch w=0.27u l=0.06u
.ends
.subckt SDFKSND0 SI D SE CP SN Q QN VDD VSS
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI49-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.15u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI141-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI142-M_u2 QN net69 VSS VSS nch w=0.195u l=0.06u
MI72-M_u2 net116 SN VSS VSS nch w=0.15u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.24u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI78 net132 net116 VSS VSS nch w=0.195u l=0.06u
MI79 net132 D VSS VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI49-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.2u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.33u l=0.06u
MI141-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI142-M_u3 QN net69 VDD VDD pch w=0.26u l=0.06u
MI72-M_u3 net116 SN VDD VDD pch w=0.2u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.51u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net116 net139 VDD pch w=0.26u l=0.06u
MI77 net139 D net132 VDD pch w=0.26u l=0.06u
.ends
.subckt SDFKSND1 SI D SE CP SN Q QN VDD VSS
MI138-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI142-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI140-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net116 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.24u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI78 net132 net116 VSS VSS nch w=0.195u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI142-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI140-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.33u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net116 SN VDD VDD pch w=0.28u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.51u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net116 net139 VDD pch w=0.28u l=0.06u
MI77 net139 D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKSND2 SI D SE CP SN Q QN VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI142-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net123 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.24u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI78 net132 net123 VSS VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.33u l=0.06u
MI142-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net123 SN VDD VDD pch w=0.28u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.51u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net123 net145 VDD pch w=0.28u l=0.06u
MI77 net145 D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKSND4 SI D SE CP SN Q QN VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI146-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI136-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI142-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.42u l=0.06u
MI115-M_u2 net69 net105 VSS VSS nch w=0.245u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI143-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI141-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI144-M_u2 QN net69 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net123 SN VSS VSS nch w=0.195u l=0.06u
MI145-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.535u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI78 net132 net123 VSS VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI146-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI136-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI142-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.68u l=0.06u
MI115-M_u3 net69 net105 VDD VDD pch w=0.33u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI143-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI141-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI144-M_u3 QN net69 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net123 SN VDD VDD pch w=0.28u l=0.06u
MI145-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net123 net145 VDD pch w=0.28u l=0.06u
MI77 net145 D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKSNQD0 SI D SE CP SN Q VDD VSS
MI64 net77 net85 VSS VSS nch w=0.195u l=0.06u
MI65 net146 net81 net77 VSS nch w=0.195u l=0.06u
MI62 net146 SE net102 VSS nch w=0.15u l=0.06u
MI89 net158 INCP net87 VSS nch w=0.15u l=0.06u
MI90 net87 net93 VSS VSS nch w=0.15u l=0.06u
MI106 net93 INCP net69 VSS nch w=0.21u l=0.06u
MI122 net068 Q VSS VSS nch w=0.15u l=0.06u
MI135 net69 INCPB net068 VSS nch w=0.15u l=0.06u
MI83 net158 INCPB net146 VSS nch w=0.23u l=0.06u
MI63 net102 net0102 VSS VSS nch w=0.15u l=0.06u
MI78 net81 net83 VSS VSS nch w=0.195u l=0.06u
MI79 net81 D VSS VSS nch w=0.195u l=0.06u
MI115-M_u2 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net85 SE VSS VSS nch w=0.15u l=0.06u
MI116-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net158 VSS VSS nch w=0.34u l=0.06u
MI109-M_u2 Q net69 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net83 SN VSS VSS nch w=0.15u l=0.06u
MI115-M_u3 net0102 SI VDD VDD pch w=0.2u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI45-M_u3 net85 SE VDD VDD pch w=0.2u l=0.06u
MI116-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net158 VDD VDD pch w=0.34u l=0.06u
MI109-M_u3 Q net69 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net83 SN VDD VDD pch w=0.2u l=0.06u
MI123 net69 INCP net0115 VDD pch w=0.15u l=0.06u
MI50 net130 SE VDD VDD pch w=0.255u l=0.06u
MI82 net158 INCP net117 VDD pch w=0.3u l=0.06u
MI53 net117 net85 net145 VDD pch w=0.15u l=0.06u
MI88 net150 net93 VDD VDD pch w=0.15u l=0.06u
MI51 net117 net81 net130 VDD pch w=0.255u l=0.06u
MI52 net145 net0102 VDD VDD pch w=0.15u l=0.06u
MI87 net158 INCPB net150 VDD pch w=0.15u l=0.06u
MI136 net0115 Q VDD VDD pch w=0.15u l=0.06u
MI113 net93 INCPB net69 VDD pch w=0.43u l=0.06u
MI75 VDD net83 net166 VDD pch w=0.26u l=0.06u
MI77 net166 D net81 VDD pch w=0.26u l=0.06u
.ends
.subckt SDFKSNQD1 SI D SE CP SN Q VDD VSS
MI142-M_u2 net69 net105 VSS VSS nch w=0.15u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI141-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI140-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net116 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.24u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI78 net132 net116 VSS VSS nch w=0.195u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI142-M_u3 net69 net105 VDD VDD pch w=0.15u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI141-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI140-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.33u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net116 SN VDD VDD pch w=0.28u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.51u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net116 net139 VDD pch w=0.28u l=0.06u
MI77 net139 D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKSNQD2 SI D SE CP SN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI142-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI141-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI144-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI72-M_u2 net123 SN VSS VSS nch w=0.195u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.24u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.26u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI78 net132 net123 VSS VSS nch w=0.195u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI142-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI141-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net93 net155 VDD VDD pch w=0.33u l=0.06u
MI144-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI72-M_u3 net123 SN VDD VDD pch w=0.26u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.51u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI75 VDD net123 net145 VDD pch w=0.28u l=0.06u
MI77 net145 D net132 VDD pch w=0.52u l=0.06u
.ends
.subckt SDFKSNQD4 SI D SE CP SN Q VDD VSS
MI138-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI130-M_u2 net109 net90 VSS VSS nch w=0.39u l=0.06u
MI145-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI146-M_u2 net107 SE VSS VSS nch w=0.195u l=0.06u
MI72-M_u2 net235 SN VSS VSS nch w=0.195u l=0.06u
MI139-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI140-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI42_0-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI42_1-M_u2 net93 net155 VSS VSS nch w=0.21u l=0.06u
MI147-M_u2 net69 net105 VSS VSS nch w=0.195u l=0.06u
MI116-M_u2 Q net105 VSS VSS nch w=0.39u l=0.06u
MI112 net93 INCP net105 VSS nch w=0.535u l=0.06u
MI135 net87 SI VSS VSS nch w=0.15u l=0.06u
MI128 net132 net107 net90 VSS nch w=0.2u l=0.06u
MI29 net105 INCPB net79 VSS nch w=0.15u l=0.06u
MI26 net79 net69 VSS VSS nch w=0.15u l=0.06u
MI126 net109 INCPB net155 VSS nch w=0.27u l=0.06u
MI101 net155 INCP net95 VSS nch w=0.15u l=0.06u
MI102 net95 net93 VSS VSS nch w=0.15u l=0.06u
MI78 net132 net235 VSS VSS nch w=0.195u l=0.06u
MI79 net132 D VSS VSS nch w=0.39u l=0.06u
MI134 net90 SE net87 VSS nch w=0.15u l=0.06u
MI138-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI130-M_u3 net109 net90 VDD VDD pch w=0.51u l=0.06u
MI145-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI146-M_u3 net107 SE VDD VDD pch w=0.26u l=0.06u
MI72-M_u3 net235 SN VDD VDD pch w=0.26u l=0.06u
MI139-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI140-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI42_0-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI42_1-M_u3 net93 net155 VDD VDD pch w=0.34u l=0.06u
MI147-M_u3 net69 net105 VDD VDD pch w=0.26u l=0.06u
MI116-M_u3 Q net105 VDD VDD pch w=0.52u l=0.06u
MI28 net105 INCP net168 VDD pch w=0.15u l=0.06u
MI129 net132 SE net90 VDD pch w=0.38u l=0.06u
MI24 net168 net69 VDD VDD pch w=0.15u l=0.06u
MI133 net138 net107 net90 VDD pch w=0.2u l=0.06u
MI119 net93 INCPB net105 VDD pch w=0.97u l=0.06u
MI127 net109 INCP net155 VDD pch w=0.34u l=0.06u
MI99 net155 INCPB net153 VDD pch w=0.15u l=0.06u
MI100 net153 net93 VDD VDD pch w=0.15u l=0.06u
MI131 VDD SI net138 VDD pch w=0.2u l=0.06u
MI77 net265 D net132 VDD pch w=0.52u l=0.06u
MI75 VDD net235 net265 VDD pch w=0.28u l=0.06u
.ends
.subckt SDFNCND0 SI D SE CPN CDN Q QN VDD VSS
MI162 net177 D net072 VSS nch w=0.26u l=0.06u
MI150 net62 net101 d2 VSS nch w=0.15u l=0.06u
MI149 d1 INCPB d2 VSS nch w=0.2u l=0.06u
MI49 net79 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net82 d1 net79 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net82 VSS nch w=0.15u l=0.06u
MI77 d0 net101 net177 VSS nch w=0.16u l=0.06u
MI78 net89 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net89 VSS nch w=0.15u l=0.06u
MI81 net072 net120 VSS VSS nch w=0.26u l=0.06u
MI167-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI168-M_u2 QN net62 VSS VSS nch w=0.195u l=0.06u
MI172-M_u2 net62 d3 VSS VSS nch w=0.195u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.15u l=0.06u
MI165-M_u2 INCPB CPN VSS VSS nch w=0.15u l=0.06u
MI171-M_u2 net101 INCPB VSS VSS nch w=0.195u l=0.06u
MI173-M_u4 XI173-net6 CDN VSS VSS nch w=0.35u l=0.06u
MI173-M_u3 d3 d2 XI173-net6 VSS nch w=0.35u l=0.06u
MI167-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI168-M_u3 QN net62 VDD VDD pch w=0.26u l=0.06u
MI172-M_u3 net62 d3 VDD VDD pch w=0.26u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.2u l=0.06u
MI165-M_u3 INCPB CPN VDD VDD pch w=0.2u l=0.06u
MI171-M_u3 net101 INCPB VDD VDD pch w=0.26u l=0.06u
MI164 net117 D net69 VDD pch w=0.33u l=0.06u
MI155 net62 INCPB d2 VDD pch w=0.15u l=0.06u
MI45 d0 net101 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI163 net117 net120 net142 VDD pch w=0.15u l=0.06u
MI73 net69 SE VDD VDD pch w=0.33u l=0.06u
MI74 d0 INCPB net117 VDD pch w=0.49u l=0.06u
MI75 net142 SI VDD VDD pch w=0.15u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 net101 d2 VDD pch w=0.29u l=0.06u
MI173-M_u2 d3 CDN VDD VDD pch w=0.44u l=0.06u
MI173-M_u1 d3 d2 VDD VDD pch w=0.44u l=0.06u
.ends
.subckt SDFNCND1 SI D SE CPN CDN Q QN VDD VSS
MI162 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI150 net62 net101 d2 VSS nch w=0.15u l=0.06u
MI149 d1 INCPB d2 VSS nch w=0.2u l=0.06u
MI49 net79 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net82 d1 net79 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net82 VSS nch w=0.15u l=0.06u
MI77 d0 net101 net177 VSS nch w=0.16u l=0.06u
MI78 net89 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net89 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.4u l=0.06u
MI151-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI179-M_u2 net62 d3 VSS VSS nch w=0.195u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.23u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI165-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI178-M_u2 net101 INCPB VSS VSS nch w=0.195u l=0.06u
MI180-M_u4 XI180-net6 CDN VSS VSS nch w=0.35u l=0.06u
MI180-M_u3 d3 d2 XI180-net6 VSS nch w=0.35u l=0.06u
MI151-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI179-M_u3 net62 d3 VDD VDD pch w=0.26u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI165-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI178-M_u3 net101 INCPB VDD VDD pch w=0.26u l=0.06u
MI164 net117 SE net69 VDD pch w=0.44u l=0.06u
MI155 net62 INCPB d2 VDD pch w=0.15u l=0.06u
MI45 d0 net101 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI163 net117 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.51u l=0.06u
MI74 d0 INCPB net117 VDD pch w=0.49u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 net101 d2 VDD pch w=0.29u l=0.06u
MI180-M_u2 d3 CDN VDD VDD pch w=0.44u l=0.06u
MI180-M_u1 d3 d2 VDD VDD pch w=0.44u l=0.06u
.ends
.subckt SDFNCND2 SI D SE CPN CDN Q QN VDD VSS
MI162 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI150 net62 net101 d2 VSS nch w=0.15u l=0.06u
MI149 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net79 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net82 d1 net79 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net82 VSS nch w=0.15u l=0.06u
MI77 d0 net101 net177 VSS nch w=0.17u l=0.06u
MI78 net89 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net89 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.4u l=0.06u
MI165-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI159-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI160-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI151-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI153-M_u2 net62 d3 VSS VSS nch w=0.23u l=0.06u
MI168-M_u2 net101 INCPB VSS VSS nch w=0.195u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI158-M_u4 XI158-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158-M_u3 d3 d2 XI158-net6 VSS nch w=0.23u l=0.06u
MI167-M_u4 XI167-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI167-M_u3 d3 d2 XI167-net6 VSS nch w=0.23u l=0.06u
MI165-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI159-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI160-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI151-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI153-M_u3 net62 d3 VDD VDD pch w=0.33u l=0.06u
MI168-M_u3 net101 INCPB VDD VDD pch w=0.26u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.34u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI164 net117 SE net69 VDD pch w=0.44u l=0.06u
MI155 net62 INCPB d2 VDD pch w=0.15u l=0.06u
MI45 d0 net101 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI163 net117 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.51u l=0.06u
MI74 d0 INCPB net117 VDD pch w=0.49u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 net101 d2 VDD pch w=0.4u l=0.06u
MI158-M_u2 d3 CDN VDD VDD pch w=0.33u l=0.06u
MI158-M_u1 d3 d2 VDD VDD pch w=0.33u l=0.06u
MI167-M_u2 d3 CDN VDD VDD pch w=0.33u l=0.06u
MI167-M_u1 d3 d2 VDD VDD pch w=0.33u l=0.06u
.ends
.subckt SDFNCND4 SI D SE CPN CDN Q QN VDD VSS
MI162 net177 net120 net69 VSS nch w=0.35u l=0.06u
MI150 net62 net101 d2 VSS nch w=0.15u l=0.06u
MI149 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net79 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net82 d1 net79 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net82 VSS nch w=0.15u l=0.06u
MI77 d0 net101 net177 VSS nch w=0.17u l=0.06u
MI78 net89 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net89 VSS nch w=0.15u l=0.06u
MI81 net69 D VSS VSS nch w=0.39u l=0.06u
MI165-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI159-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI160-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI151-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI152-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI153-M_u2 net62 d3 VSS VSS nch w=0.62u l=0.06u
MI166-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI174-M_u2 net101 INCPB VSS VSS nch w=0.39u l=0.06u
MI167-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI168-M_u2 QN net62 VSS VSS nch w=0.39u l=0.06u
MI85-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI173-M_u2 INCPB CPN VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI158-M_u4 XI158-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI158-M_u3 d3 d2 XI158-net6 VSS nch w=0.23u l=0.06u
MI170-M_u4 XI170-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI170-M_u3 d3 d2 XI170-net6 VSS nch w=0.23u l=0.06u
MI165-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI159-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI160-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI151-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI153-M_u3 net62 d3 VDD VDD pch w=0.85u l=0.06u
MI166-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI174-M_u3 net101 INCPB VDD VDD pch w=0.52u l=0.06u
MI167-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI168-M_u3 QN net62 VDD VDD pch w=0.52u l=0.06u
MI85-M_u3 d1 d0 VDD VDD pch w=0.34u l=0.06u
MI173-M_u3 INCPB CPN VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI164 net117 SE net69 VDD pch w=0.44u l=0.06u
MI155 net62 INCPB d2 VDD pch w=0.15u l=0.06u
MI45 d0 net101 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI163 net117 net120 net142 VDD pch w=0.2u l=0.06u
MI73 net69 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net117 VDD pch w=0.47u l=0.06u
MI75 net142 SI VDD VDD pch w=0.2u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI154 d1 net101 d2 VDD pch w=0.4u l=0.06u
MI158-M_u2 d3 CDN VDD VDD pch w=0.33u l=0.06u
MI158-M_u1 d3 d2 VDD VDD pch w=0.33u l=0.06u
MI170-M_u2 d3 CDN VDD VDD pch w=0.33u l=0.06u
MI170-M_u1 d3 d2 VDD VDD pch w=0.33u l=0.06u
.ends
.subckt SDFNCSND0 SI D SE CPN CDN SDN Q QN VDD VSS
MI91 d4 net105 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net86 VSS nch w=0.15u l=0.06u
MI77 d0 net105 net177 VSS nch w=0.17u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI79 net96 net120 VSS VSS nch w=0.26u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net177 D net96 VSS nch w=0.26u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.15u l=0.06u
MI31-M_u2 INCPB CPN VSS VSS nch w=0.15u l=0.06u
MI100-M_u2 net105 INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.15u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.15u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.2u l=0.06u
MI31-M_u3 INCPB CPN VDD VDD pch w=0.2u l=0.06u
MI100-M_u3 net105 INCPB VDD VDD pch w=0.26u l=0.06u
MI45 d0 net105 net166 VDD pch w=0.15u l=0.06u
MI43 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.15u l=0.06u
MI72 net149 SE VDD VDD pch w=0.33u l=0.06u
MI73 net104 D net149 VDD pch w=0.33u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.49u l=0.06u
MI75 net148 SI VDD VDD pch w=0.15u l=0.06u
MI98 d1 net105 d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.2u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFNCSND1 SI D SE CPN CDN SDN Q QN VDD VSS
MI91 d4 net105 d2 VSS nch w=0.15u l=0.06u
MI102 net177 net120 net84 VSS nch w=0.35u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net86 VSS nch w=0.15u l=0.06u
MI77 d0 net105 net177 VSS nch w=0.17u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net84 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI108-M_u2 net105 INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI103-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI108-M_u3 net105 INCPB VDD VDD pch w=0.26u l=0.06u
MI101 net104 SE net84 VDD pch w=0.44u l=0.06u
MI105 d0 net105 net166 VDD pch w=0.15u l=0.06u
MI104 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net84 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.49u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 net105 d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFNCSND2 SI D SE CPN CDN SDN Q QN VDD VSS
MI91 d4 net105 d2 VSS nch w=0.15u l=0.06u
MI102 net177 net120 net84 VSS nch w=0.35u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net86 VSS nch w=0.15u l=0.06u
MI77 d0 net105 net177 VSS nch w=0.17u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net84 D VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI100-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI104-M_u2 net105 INCPB VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI100-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI104-M_u3 net105 INCPB VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI101 net104 SE net84 VDD pch w=0.44u l=0.06u
MI107 d0 net105 net166 VDD pch w=0.15u l=0.06u
MI106 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net84 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.49u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 net105 d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.38u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.38u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFNCSND4 SI D SE CPN CDN SDN Q QN VDD VSS
MI91 d4 net105 d2 VSS nch w=0.15u l=0.06u
MI102 net177 net120 net84 VSS nch w=0.35u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.19u l=0.06u
MI49 net83 CDN VSS VSS nch w=0.15u l=0.06u
MI48 net86 d1 net83 VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net86 VSS nch w=0.15u l=0.06u
MI77 d0 net105 net177 VSS nch w=0.17u l=0.06u
MI78 net93 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net93 VSS nch w=0.15u l=0.06u
MI81 net84 D VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI95-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI96-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI100-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI104-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI105-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI114-M_u2 INCPB CPN VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI115-M_u2 net105 INCPB VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.35u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.35u l=0.06u
MI94-M_u4 XI94-net6 d2 VSS VSS nch w=0.17u l=0.06u
MI94-M_u3 d3 CDN XI94-net6 VSS nch w=0.17u l=0.06u
MI107-M_u4 XI107-net6 d2 VSS VSS nch w=0.35u l=0.06u
MI107-M_u3 d3 CDN XI107-net6 VSS nch w=0.35u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.21u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.21u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI95-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI96-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI100-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI104-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI105-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI114-M_u3 INCPB CPN VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI115-M_u3 net105 INCPB VDD VDD pch w=0.52u l=0.06u
MI101 net104 SE net84 VDD pch w=0.44u l=0.06u
MI109 d0 net105 net166 VDD pch w=0.15u l=0.06u
MI108 net166 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net148 VDD pch w=0.2u l=0.06u
MI73 net84 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.45u l=0.06u
MI75 net148 SI VDD VDD pch w=0.2u l=0.06u
MI98 d1 net105 d2 VDD pch w=0.32u l=0.06u
MI44 net166 CDN VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.38u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.38u l=0.06u
MI94-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI94-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI107-M_u2 d3 d2 VDD VDD pch w=0.32u l=0.06u
MI107-M_u1 d3 CDN VDD VDD pch w=0.32u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.4u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SDFND0 SI D SE CPN Q QN VDD VSS
MI25 net65 INCPB d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCPB net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 net89 d2 VSS nch w=0.15u l=0.06u
MU65 net28 net89 net37 VSS nch w=0.21u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU64 net81 net57 VSS VSS nch w=0.26u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net37 D net81 VSS nch w=0.26u l=0.06u
MI39-M_u2 net55 d3 VSS VSS nch w=0.15u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.195u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.15u l=0.06u
MU84-M_u2 INCPB CPN VSS VSS nch w=0.15u l=0.06u
MI38-M_u2 net89 INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI39-M_u3 net55 d3 VDD VDD pch w=0.2u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.26u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.2u l=0.06u
MU84-M_u3 INCPB CPN VDD VDD pch w=0.2u l=0.06u
MI38-M_u3 net89 INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCPB d2 VDD pch w=0.15u l=0.06u
MI36 net65 net89 d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.15u l=0.06u
MU60 net128 SE VDD VDD pch w=0.33u l=0.06u
MU61 net13 D net128 VDD pch w=0.33u l=0.06u
MU62 net28 INCPB net13 VDD pch w=0.28u l=0.06u
MU70 net132 SI VDD VDD pch w=0.15u l=0.06u
MI10 net28 net89 net137 VDD pch w=0.15u l=0.06u
.ends
.subckt SDFND1 SI D SE CPN Q QN VDD VSS
MI39 net37 net57 net110 VSS nch w=0.35u l=0.06u
MI25 net65 INCPB d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCPB net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 net89 d2 VSS nch w=0.15u l=0.06u
MU65 net28 net89 net37 VSS nch w=0.21u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net110 D VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.195u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MI41-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI43-M_u2 net89 INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=0.26u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MI41-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI43-M_u3 net89 INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCPB d2 VDD pch w=0.15u l=0.06u
MI40 net13 SE net110 VDD pch w=0.44u l=0.06u
MI36 net65 net89 d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net110 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCPB net13 VDD pch w=0.28u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 net89 net137 VDD pch w=0.15u l=0.06u
.ends
.subckt SDFND2 SI D SE CPN Q QN VDD VSS
MI39 net37 net57 net110 VSS nch w=0.35u l=0.06u
MI25 net65 INCPB d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCPB net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 net89 d2 VSS nch w=0.15u l=0.06u
MU65 net28 net89 net37 VSS nch w=0.21u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net110 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI38-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI41-M_u2 net89 INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI38-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI41-M_u3 net89 INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCPB d2 VDD pch w=0.15u l=0.06u
MI40 net13 SE net110 VDD pch w=0.44u l=0.06u
MI36 net65 net89 d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net110 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCPB net13 VDD pch w=0.28u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 net89 net137 VDD pch w=0.15u l=0.06u
.ends
.subckt SDFND4 SI D SE CPN Q QN VDD VSS
MI39 net37 net57 net110 VSS nch w=0.35u l=0.06u
MI25 net65 INCPB d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCPB net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI26 net55 net89 d2 VSS nch w=0.15u l=0.06u
MU65 net28 net89 net37 VSS nch w=0.21u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net110 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI38-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI28-M_u2 net55 d3 VSS VSS nch w=0.78u l=0.06u
MI30_0-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI30_1-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI41-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI43-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI44-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI34-M_u2 QN net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CPN VSS VSS nch w=0.39u l=0.06u
MU85-M_u2 net89 INCPB VSS VSS nch w=0.39u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI38-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI28-M_u3 net55 d3 VDD VDD pch w=1.04u l=0.06u
MI30_0-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI30_1-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI41-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI43-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI44-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI34-M_u3 QN net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CPN VDD VDD pch w=0.52u l=0.06u
MU85-M_u3 net89 INCPB VDD VDD pch w=0.52u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI35 net55 INCPB d2 VDD pch w=0.15u l=0.06u
MI40 net13 SE net110 VDD pch w=0.44u l=0.06u
MI36 net65 net89 d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net110 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCPB net13 VDD pch w=0.28u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 net89 net137 VDD pch w=0.15u l=0.06u
.ends
.subckt SDFNSND0 SI D SE CPN SDN Q QN VDD VSS
MI91 d4 net95 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.39u l=0.06u
MI101 net177 D net76 VSS nch w=0.26u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net72 VSS nch w=0.15u l=0.06u
MI77 d0 net95 net177 VSS nch w=0.17u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net76 net095 VSS VSS nch w=0.26u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net095 SE VSS VSS nch w=0.15u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CPN VSS VSS nch w=0.15u l=0.06u
MI105-M_u2 net95 INCPB VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 QN d4 VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.15u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.15u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net095 SE VDD VDD pch w=0.2u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CPN VDD VDD pch w=0.2u l=0.06u
MI105-M_u3 net95 INCPB VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 QN d4 VDD VDD pch w=0.26u l=0.06u
MI102 net104 D net0117 VDD pch w=0.33u l=0.06u
MI45 d0 net95 net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net095 net131 VDD pch w=0.15u l=0.06u
MI73 net0117 SE VDD VDD pch w=0.33u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.47u l=0.06u
MI75 net131 SI VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI98 d1 net95 d2 VDD pch w=0.315u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFNSND1 SI D SE CPN SDN Q QN VDD VSS
MI91 d4 net95 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.39u l=0.06u
MI101 net177 net120 net76 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net72 VSS nch w=0.15u l=0.06u
MI77 d0 net95 net177 VSS nch w=0.17u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net76 D VSS VSS nch w=0.39u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI104-M_u2 net95 INCPB VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI104-M_u3 net95 INCPB VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI102 net104 SE net76 VDD pch w=0.44u l=0.06u
MI45 d0 net95 net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net76 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.49u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI98 d1 net95 d2 VDD pch w=0.315u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFNSND2 SI D SE CPN SDN Q QN VDD VSS
MI91 d4 net95 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.39u l=0.06u
MI101 net177 net120 net76 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net72 VSS nch w=0.15u l=0.06u
MI77 d0 net95 net177 VSS nch w=0.17u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net76 D VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 net95 INCPB VSS VSS nch w=0.195u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI100-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI104-M_u2 INCPB CPN VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI95-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.39u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.39u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI103-M_u3 net95 INCPB VDD VDD pch w=0.26u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI100-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI104-M_u3 INCPB CPN VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI95-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI102 net104 SE net76 VDD pch w=0.44u l=0.06u
MI45 d0 net95 net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net76 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.47u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI98 d1 net95 d2 VDD pch w=0.315u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.52u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.52u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFNSND4 SI D SE CPN SDN Q QN VDD VSS
MI91 d4 net95 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCPB d2 VSS nch w=0.39u l=0.06u
MI101 net177 net120 net76 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCPB net72 VSS nch w=0.15u l=0.06u
MI77 d0 net95 net177 VSS nch w=0.17u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net76 D VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI110-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI109-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI111-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI114-M_u2 INCPB CPN VSS VSS nch w=0.39u l=0.06u
MI107-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI112-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96_0-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI96_1-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI115-M_u2 net95 INCPB VSS VSS nch w=0.39u l=0.06u
MI113-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.39u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.39u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI108-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI110-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI109-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI111-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI114-M_u3 INCPB CPN VDD VDD pch w=0.52u l=0.06u
MI107-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI112-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96_0-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI96_1-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI115-M_u3 net95 INCPB VDD VDD pch w=0.52u l=0.06u
MI113-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI102 net104 SE net76 VDD pch w=0.44u l=0.06u
MI45 d0 net95 net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net76 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCPB net104 VDD pch w=0.47u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI97 d4 INCPB d2 VDD pch w=0.15u l=0.06u
MI98 d1 net95 d2 VDD pch w=0.315u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.52u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.52u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFQD0 SI D SE CP Q VDD VSS
MI39 net117 d3 VSS VSS nch w=0.15u l=0.06u
MI29 d2 INCPB net117 VSS nch w=0.15u l=0.06u
MI25 net110 INCP d2 VSS nch w=0.15u l=0.06u
MI13 net69 INCP net109 VSS nch w=0.15u l=0.06u
MI14 net109 net110 VSS VSS nch w=0.15u l=0.06u
MU65 net69 INCPB net97 VSS nch w=0.15u l=0.06u
MU67 net103 SI VSS VSS nch w=0.15u l=0.06u
MI51 net97 net78 VSS VSS nch w=0.15u l=0.06u
MI42 net78 D net94 VSS nch w=0.23u l=0.06u
MU68 net78 SE net103 VSS nch w=0.15u l=0.06u
MU63 net94 net131 VSS VSS nch w=0.23u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.15u l=0.06u
MI49-M_u2 Q d2 VSS VSS nch w=0.15u l=0.06u
MU71-M_u2 net131 SE VSS VSS nch w=0.19u l=0.06u
MI43-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI46-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net110 net69 VSS VSS nch w=0.21u l=0.06u
MI24 net87 d3 VDD VDD pch w=0.15u l=0.06u
MI11 net65 net110 VDD VDD pch w=0.15u l=0.06u
MI50 net057 net78 VDD VDD pch w=0.25u l=0.06u
MI36 net110 INCPB d2 VDD pch w=0.35u l=0.06u
MU69 net78 net131 net80 VDD pch w=0.15u l=0.06u
MI41 net78 D net77 VDD pch w=0.3u l=0.06u
MU61 net77 SE VDD VDD pch w=0.38u l=0.06u
MU62 net69 INCP net057 VDD pch w=0.25u l=0.06u
MU70 net80 SI VDD VDD pch w=0.15u l=0.06u
MI10 net69 INCPB net65 VDD pch w=0.15u l=0.06u
MI38 d2 INCP net87 VDD pch w=0.15u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.15u l=0.06u
MI49-M_u3 Q d2 VDD VDD pch w=0.24u l=0.06u
MU71-M_u3 net131 SE VDD VDD pch w=0.26u l=0.06u
MI43-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI46-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net110 net69 VDD VDD pch w=0.335u l=0.06u
.ends
.subckt SDFQD1 SI D SE CP Q VDD VSS
MI30-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MI43-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI46-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI39 net60 d3 VSS VSS nch w=0.15u l=0.06u
MI29 d2 INCPB net60 VSS nch w=0.15u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.18u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MI42 net37 net57 net13 VSS nch w=0.35u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net13 D VSS VSS nch w=0.39u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MI43-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI46-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI38 d2 INCP net62 VDD pch w=0.15u l=0.06u
MI24 net62 d3 VDD VDD pch w=0.15u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net120 net57 net132 VDD pch w=0.2u l=0.06u
MI41 net120 SE net13 VDD pch w=0.44u l=0.06u
MU61 net13 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net120 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
.ends
.subckt SDFQD2 SI D SE CP Q VDD VSS
MI39 net37 net57 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI45 net061 d3 VSS VSS nch w=0.15u l=0.06u
MI29 d2 INCPB net061 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.15u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI46-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI33-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI46-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI33-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI24 net0110 d3 VDD VDD pch w=0.15u l=0.06u
MI38 d2 INCP net0110 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFQD4 SI D SE CP Q VDD VSS
MI39 net37 net57 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI29 d2 INCPB net0155 VSS nch w=0.15u l=0.06u
MI49 net0155 net55 VSS VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.17u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI37-M_u2 Q net55 VSS VSS nch w=0.39u l=0.06u
MI50-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI51-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI44-M_u2 Q net55 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 net55 d2 VSS VSS nch w=0.78u l=0.06u
MI45-M_u2 Q net55 VSS VSS nch w=0.39u l=0.06u
MI33-M_u2 Q net55 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI37-M_u3 Q net55 VDD VDD pch w=0.52u l=0.06u
MI50-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI51-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI44-M_u3 Q net55 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 net55 d2 VDD VDD pch w=1.04u l=0.06u
MI45-M_u3 Q net55 VDD VDD pch w=0.52u l=0.06u
MI33-M_u3 Q net55 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI38 d2 INCP net0203 VDD pch w=0.15u l=0.06u
MI24 net0203 net55 VDD VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.3u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFQND0 SI D SE CP QN VDD VSS
MI30-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.15u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI44-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI39 net37 D net64 VSS nch w=0.26u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI41 net054 QN VSS VSS nch w=0.15u l=0.06u
MI29 d2 INCPB net054 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.16u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 net57 VSS VSS nch w=0.26u l=0.06u
MI30-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.2u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI44-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI24 net064 QN VDD VDD pch w=0.15u l=0.06u
MI38 d2 INCP net064 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.15u l=0.06u
MU61 net0111 SE VDD VDD pch w=0.33u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.33u l=0.06u
MU70 net132 SI VDD VDD pch w=0.15u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 D net0111 VDD pch w=0.33u l=0.06u
.ends
.subckt SDFQND1 SI D SE CP QN VDD VSS
MI39 net37 net57 net64 VSS nch w=0.35u l=0.06u
MI25 net65 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net28 INCP net66 VSS nch w=0.15u l=0.06u
MI14 net66 net65 VSS VSS nch w=0.15u l=0.06u
MI45 net054 net55 VSS VSS nch w=0.15u l=0.06u
MI44 d2 INCPB net054 VSS nch w=0.15u l=0.06u
MU65 net28 INCPB net37 VSS nch w=0.16u l=0.06u
MU67 net83 SI VSS VSS nch w=0.15u l=0.06u
MU68 net37 SE net83 VSS nch w=0.15u l=0.06u
MU63 net64 D VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 net55 d2 VSS VSS nch w=0.15u l=0.06u
MI49-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net57 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net65 net28 VSS VSS nch w=0.35u l=0.06u
MI30-M_u3 net55 d2 VDD VDD pch w=0.15u l=0.06u
MI49-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net57 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net65 net28 VDD VDD pch w=0.38u l=0.06u
MI11 net137 net65 VDD VDD pch w=0.15u l=0.06u
MI46 net098 net55 VDD VDD pch w=0.15u l=0.06u
MI47 d2 INCP net098 VDD pch w=0.15u l=0.06u
MI36 net65 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net13 net57 net132 VDD pch w=0.2u l=0.06u
MU61 net64 D VDD VDD pch w=0.52u l=0.06u
MU62 net28 INCP net13 VDD pch w=0.33u l=0.06u
MU70 net132 SI VDD VDD pch w=0.2u l=0.06u
MI10 net28 INCPB net137 VDD pch w=0.15u l=0.06u
MI40 net13 SE net64 VDD pch w=0.44u l=0.06u
.ends
.subckt SDFQND2 SI D SE CP QN VDD VSS
MI11 net83 net120 VDD VDD pch w=0.15u l=0.06u
MI46 net79 net98 VDD VDD pch w=0.15u l=0.06u
MI47 d2 INCP net79 VDD pch w=0.15u l=0.06u
MI40 net71 SE net101 VDD pch w=0.44u l=0.06u
MI36 net120 INCPB d2 VDD pch w=0.44u l=0.06u
MU69 net71 net94 net73 VDD pch w=0.2u l=0.06u
MU61 net101 D VDD VDD pch w=0.52u l=0.06u
MU62 net65 INCP net71 VDD pch w=0.33u l=0.06u
MU70 net73 SI VDD VDD pch w=0.2u l=0.06u
MI10 net65 INCPB net83 VDD pch w=0.15u l=0.06u
MI30-M_u3 net98 d2 VDD VDD pch w=0.15u l=0.06u
MI49-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net94 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI50-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU72-M_u3 net120 net65 VDD VDD pch w=0.38u l=0.06u
MI30-M_u2 net98 d2 VSS VSS nch w=0.15u l=0.06u
MI49-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net94 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI50-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU72-M_u2 net120 net65 VSS VSS nch w=0.35u l=0.06u
MU68 net104 SE net103 VSS nch w=0.15u l=0.06u
MI39 net104 net94 net101 VSS nch w=0.35u l=0.06u
MU63 net101 D VSS VSS nch w=0.39u l=0.06u
MI25 net120 INCP d2 VSS nch w=0.22u l=0.06u
MI13 net65 INCP net119 VSS nch w=0.15u l=0.06u
MI14 net119 net120 VSS VSS nch w=0.15u l=0.06u
MI45 net112 net98 VSS VSS nch w=0.15u l=0.06u
MI44 d2 INCPB net112 VSS nch w=0.15u l=0.06u
MU65 net65 INCPB net104 VSS nch w=0.16u l=0.06u
MU67 net103 SI VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SDFQND4 SI D SE CP QN VDD VSS
MI13 net66 INCP net77 VSS nch w=0.15u l=0.06u
MI14 net77 net76 VSS VSS nch w=0.15u l=0.06u
MI25 net76 INCP d2 VSS nch w=0.22u l=0.06u
MI44 d2 INCPB net72 VSS nch w=0.15u l=0.06u
MU67 net63 SI VSS VSS nch w=0.15u l=0.06u
MI45 net72 net110 VSS VSS nch w=0.15u l=0.06u
MU65 net66 INCPB net90 VSS nch w=0.16u l=0.06u
MU63 net84 D VSS VSS nch w=0.39u l=0.06u
MU68 net90 SE net63 VSS nch w=0.15u l=0.06u
MI39 net90 net106 net84 VSS nch w=0.35u l=0.06u
MI54-M_u2 net76 net66 VSS VSS nch w=0.35u l=0.06u
MI51-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MI52-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MI30-M_u2 net110 d2 VSS VSS nch w=0.15u l=0.06u
MI49-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MU71-M_u2 net106 SE VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI50-M_u2 QN d2 VSS VSS nch w=0.39u l=0.06u
MI42-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI54-M_u3 net76 net66 VDD VDD pch w=0.38u l=0.06u
MI51-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MI52-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MI30-M_u3 net110 d2 VDD VDD pch w=0.15u l=0.06u
MI49-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MU71-M_u3 net106 SE VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI50-M_u3 QN d2 VDD VDD pch w=0.52u l=0.06u
MI42-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI11 net139 net76 VDD VDD pch w=0.15u l=0.06u
MI46 net136 net110 VDD VDD pch w=0.15u l=0.06u
MI47 d2 INCP net136 VDD pch w=0.15u l=0.06u
MI40 net124 SE net84 VDD pch w=0.44u l=0.06u
MI36 net76 INCPB d2 VDD pch w=0.44u l=0.06u
MU70 net126 SI VDD VDD pch w=0.2u l=0.06u
MI10 net66 INCPB net139 VDD pch w=0.15u l=0.06u
MU69 net124 net106 net126 VDD pch w=0.2u l=0.06u
MU61 net84 D VDD VDD pch w=0.52u l=0.06u
MU62 net66 INCP net124 VDD pch w=0.33u l=0.06u
.ends
.subckt SDFSND0 SI D SE CP SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI79 net82 net120 VSS VSS nch w=0.26u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net177 D net82 VSS nch w=0.26u l=0.06u
MI100-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.15u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI31-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI95-M_u2 QN d4 VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.15u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.15u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI100-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.2u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI31-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI95-M_u3 QN d4 VDD VDD pch w=0.26u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI101 net104 net120 net131 VDD pch w=0.15u l=0.06u
MI72 net132 SE VDD VDD pch w=0.33u l=0.06u
MI73 net104 D net132 VDD pch w=0.33u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.15u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSND1 SI D SE CP SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI105-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI95-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI105-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI95-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSND2 SI D SE CP SDN Q QN VDD VSS
MI91 d4 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.22u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI105-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI108-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI107-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.195u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.195u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI105-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI108-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI107-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.26u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.26u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSND4 SI D SE CP SDN Q QN VDD VSS
MI91 d4 net0110 d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.22u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 net0110 net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI105-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI118-M_u2 INCP net0110 VSS VSS nch w=0.39u l=0.06u
MI107-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI109-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI117-M_u2 net0110 CP VSS VSS nch w=0.39u l=0.06u
MI110-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI111-M_u2 QN d4 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.39u l=0.06u
MI93-M_u3 d4 SDN XI93-net6 VSS nch w=0.39u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI105-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI118-M_u3 INCP net0110 VDD VDD pch w=0.52u l=0.06u
MI107-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI108-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI109-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI117-M_u3 net0110 CP VDD VDD pch w=0.52u l=0.06u
MI110-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI111-M_u3 QN d4 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI45 d0 net0110 net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 d4 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 net0110 d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 d4 d3 VDD VDD pch w=0.52u l=0.06u
MI93-M_u1 d4 SDN VDD VDD pch w=0.52u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSNQD0 SI D SE CP SDN Q VDD VSS
MI91 net64 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI79 net82 net120 VSS VSS nch w=0.26u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net177 D net82 VSS nch w=0.26u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.15u l=0.06u
MI101-M_u2 d3 d2 VSS VSS nch w=0.195u l=0.06u
MI31-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI100-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.2u l=0.06u
MI93-M_u3 net64 SDN XI93-net6 VSS nch w=0.2u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.2u l=0.06u
MI101-M_u3 d3 d2 VDD VDD pch w=0.26u l=0.06u
MI31-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI100-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.15u l=0.06u
MI72 net132 SE VDD VDD pch w=0.33u l=0.06u
MI73 net104 D net132 VDD pch w=0.33u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.15u l=0.06u
MI97 net64 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 net64 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 net64 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSNQD1 SI D SE CP SDN Q VDD VSS
MI91 net068 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI106-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.2u l=0.06u
MI93-M_u3 net068 SDN XI93-net6 VSS nch w=0.2u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI106-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI105 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 net068 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 net068 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 net068 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSNQD2 SI D SE CP SDN Q VDD VSS
MI91 net075 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI99-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI94-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI105-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96-M_u2 d3 d2 VSS VSS nch w=0.78u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.2u l=0.06u
MI93-M_u3 net075 SDN XI93-net6 VSS nch w=0.2u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI99-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI94-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI105-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96-M_u3 d3 d2 VDD VDD pch w=1.04u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 net075 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 net075 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 net075 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFSNQD4 SI D SE CP SDN Q VDD VSS
MI91 net087 INCPB d2 VSS nch w=0.15u l=0.06u
MI92 d1 INCP d2 VSS nch w=0.39u l=0.06u
MI102 net177 net120 net75 VSS nch w=0.35u l=0.06u
MI48 net72 d1 VSS VSS nch w=0.15u l=0.06u
MI47 d0 INCP net72 VSS nch w=0.15u l=0.06u
MI77 d0 INCPB net177 VSS nch w=0.24u l=0.06u
MI78 net79 SI VSS VSS nch w=0.15u l=0.06u
MI80 net177 SE net79 VSS nch w=0.15u l=0.06u
MI81 net75 D VSS VSS nch w=0.39u l=0.06u
MI108-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI109-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI111-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI103-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI107-M_u2 Q d3 VSS VSS nch w=0.39u l=0.06u
MI82-M_u2 net120 SE VSS VSS nch w=0.195u l=0.06u
MI96_0-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI96_1-M_u2 d3 d2 VSS VSS nch w=0.39u l=0.06u
MI112-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI93-M_u4 XI93-net6 d3 VSS VSS nch w=0.2u l=0.06u
MI93-M_u3 net087 SDN XI93-net6 VSS nch w=0.2u l=0.06u
MI16-M_u4 XI16-net6 d0 VSS VSS nch w=0.39u l=0.06u
MI16-M_u3 d1 SDN XI16-net6 VSS nch w=0.39u l=0.06u
MI108-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI109-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI111-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI103-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI107-M_u3 Q d3 VDD VDD pch w=0.52u l=0.06u
MI82-M_u3 net120 SE VDD VDD pch w=0.26u l=0.06u
MI96_0-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI96_1-M_u3 d3 d2 VDD VDD pch w=0.52u l=0.06u
MI112-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI45 d0 INCPB net126 VDD pch w=0.15u l=0.06u
MI43 net126 d1 VDD VDD pch w=0.15u l=0.06u
MI71 net104 net120 net131 VDD pch w=0.2u l=0.06u
MI73 net75 D VDD VDD pch w=0.52u l=0.06u
MI74 d0 INCP net104 VDD pch w=0.29u l=0.06u
MI75 net131 SI VDD VDD pch w=0.2u l=0.06u
MI101 net104 SE net75 VDD pch w=0.44u l=0.06u
MI97 net087 INCP d2 VDD pch w=0.15u l=0.06u
MI98 d1 INCPB d2 VDD pch w=0.31u l=0.06u
MI93-M_u2 net087 d3 VDD VDD pch w=0.2u l=0.06u
MI93-M_u1 net087 SDN VDD VDD pch w=0.2u l=0.06u
MI16-M_u2 d1 d0 VDD VDD pch w=0.52u l=0.06u
MI16-M_u1 d1 SDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SDFXD0 DA DB SA SI SE CP Q QN VDD VSS
MI24 net76 net72 VDD VDD pch w=0.15u l=0.06u
MI38 net138 INCP net76 VDD pch w=0.15u l=0.06u
MI153 d0 INCP net88 VDD pch w=0.3u l=0.06u
MI222 net111 net169 VDD VDD pch w=0.27u l=0.06u
MI150 net88 DA net94 VDD pch w=0.35u l=0.06u
MI233 net88 SA net91 VDD pch w=0.2u l=0.06u
MI151 net94 net128 net93 VDD pch w=0.35u l=0.06u
MI232 net91 DB net93 VDD pch w=0.2u l=0.06u
MI234 net88 net118 net90 VDD pch w=0.15u l=0.06u
MI231 net93 SE VDD VDD pch w=0.35u l=0.06u
MI235 net90 SI VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net117 VDD pch w=0.15u l=0.06u
MI102 net117 net169 VDD VDD pch w=0.15u l=0.06u
MI223 net138 INCPB net111 VDD pch w=0.27u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI229-M_u3 net128 SA VDD VDD pch w=0.2u l=0.06u
MI218-M_u3 QN net72 VDD VDD pch w=0.26u l=0.06u
MI214-M_u3 net72 net138 VDD VDD pch w=0.2u l=0.06u
MI123-M_u3 net169 d0 VDD VDD pch w=0.26u l=0.06u
MI228-M_u3 Q net138 VDD VDD pch w=0.26u l=0.06u
MI230-M_u3 net118 SE VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI41 net73 net72 VSS VSS nch w=0.15u l=0.06u
MI29 net138 INCPB net73 VSS nch w=0.15u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI229-M_u2 net128 SA VSS VSS nch w=0.15u l=0.06u
MI218-M_u2 QN net72 VSS VSS nch w=0.195u l=0.06u
MI214-M_u2 net72 net138 VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 net169 d0 VSS VSS nch w=0.195u l=0.06u
MI228-M_u2 Q net138 VSS VSS nch w=0.195u l=0.06u
MI230-M_u2 net118 SE VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI119 net158 net169 VSS VSS nch w=0.15u l=0.06u
MI240 net155 net118 VSS VSS nch w=0.355u l=0.06u
MI236 net152 SI VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net158 VSS nch w=0.15u l=0.06u
MI239 net146 DB net155 VSS nch w=0.175u l=0.06u
MI237 net153 SE net152 VSS nch w=0.15u l=0.06u
MI163 net143 SA net155 VSS nch w=0.175u l=0.06u
MI238 net153 net128 net146 VSS nch w=0.175u l=0.06u
MI160 net153 DA net143 VSS nch w=0.175u l=0.06u
MI225 net141 net169 VSS VSS nch w=0.205u l=0.06u
MI227 net138 INCP net141 VSS nch w=0.22u l=0.06u
MI164 d0 INCPB net153 VSS nch w=0.195u l=0.06u
.ends
.subckt SDFXD1 DA DB SA SI SE CP Q QN VDD VSS
MI218-M_u3 QN net098 VDD VDD pch w=0.52u l=0.06u
MI241-M_u3 net0124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0122 SA VDD VDD pch w=0.26u l=0.06u
MI228-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI214-M_u3 net098 net82 VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 net086 d0 VDD VDD pch w=0.26u l=0.06u
MI231 net0147 SE VDD VDD pch w=0.35u l=0.06u
MI233 net208 SA net0145 VDD pch w=0.435u l=0.06u
MI232 net0145 DB net0147 VDD pch w=0.255u l=0.06u
MI102 net144 net086 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net144 VDD pch w=0.15u l=0.06u
MI223 net82 INCPB net0171 VDD pch w=0.27u l=0.06u
MI234 net208 net0124 net0148 VDD pch w=0.2u l=0.06u
MI235 net0148 SI VDD VDD pch w=0.2u l=0.06u
MI222 net0171 net086 VDD VDD pch w=0.27u l=0.06u
MI150 net208 DA net162 VDD pch w=0.35u l=0.06u
MI151 net162 net0122 net0147 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net208 VDD pch w=0.3u l=0.06u
MI38 net82 INCP net070 VDD pch w=0.15u l=0.06u
MI24 net070 net098 VDD VDD pch w=0.15u l=0.06u
MI237 net265 SE net099 VSS nch w=0.15u l=0.06u
MI238 net265 net0122 net096 VSS nch w=0.175u l=0.06u
MI239 net096 DB net093 VSS nch w=0.175u l=0.06u
MI227 net82 INCP net0118 VSS nch w=0.22u l=0.06u
MI240 net093 net0124 VSS VSS nch w=0.355u l=0.06u
MI119 net79 net086 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net79 VSS nch w=0.15u l=0.06u
MI225 net0118 net086 VSS VSS nch w=0.205u l=0.06u
MI236 net099 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net265 VSS nch w=0.195u l=0.06u
MI163 net109 SA net093 VSS nch w=0.175u l=0.06u
MI160 net265 DA net109 VSS nch w=0.175u l=0.06u
MI218-M_u2 QN net098 VSS VSS nch w=0.39u l=0.06u
MI241-M_u2 net0124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0122 SA VSS VSS nch w=0.195u l=0.06u
MI228-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI214-M_u2 net098 net82 VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 net086 d0 VSS VSS nch w=0.195u l=0.06u
MI29 net82 INCPB net074 VSS nch w=0.15u l=0.06u
MI41 net074 net098 VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SDFXD2 DA DB SA SI SE CP Q QN VDD VSS
MI218-M_u3 QN net098 VDD VDD pch w=1.04u l=0.06u
MI241-M_u3 Q net82 VDD VDD pch w=1.04u l=0.06u
MI243-M_u3 net0124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0122 SA VDD VDD pch w=0.26u l=0.06u
MI214-M_u3 net098 net82 VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 net086 d0 VDD VDD pch w=0.26u l=0.06u
MI231 net0147 SE VDD VDD pch w=0.35u l=0.06u
MI233 net208 SA net0145 VDD pch w=0.435u l=0.06u
MI232 net0145 DB net0147 VDD pch w=0.255u l=0.06u
MI102 net144 net086 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net144 VDD pch w=0.15u l=0.06u
MI223 net82 INCPB net0171 VDD pch w=0.27u l=0.06u
MI234 net208 net0124 net0148 VDD pch w=0.2u l=0.06u
MI235 net0148 SI VDD VDD pch w=0.2u l=0.06u
MI222 net0171 net086 VDD VDD pch w=0.27u l=0.06u
MI150 net208 DA net162 VDD pch w=0.35u l=0.06u
MI151 net162 net0122 net0147 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net208 VDD pch w=0.3u l=0.06u
MI38 net82 INCP net070 VDD pch w=0.15u l=0.06u
MI24 net070 net098 VDD VDD pch w=0.15u l=0.06u
MI237 net265 SE net099 VSS nch w=0.15u l=0.06u
MI238 net265 net0122 net096 VSS nch w=0.175u l=0.06u
MI239 net096 DB net093 VSS nch w=0.175u l=0.06u
MI227 net82 INCP net0118 VSS nch w=0.22u l=0.06u
MI240 net093 net0124 VSS VSS nch w=0.355u l=0.06u
MI119 net79 net086 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net79 VSS nch w=0.15u l=0.06u
MI225 net0118 net086 VSS VSS nch w=0.205u l=0.06u
MI236 net099 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net265 VSS nch w=0.195u l=0.06u
MI163 net109 SA net093 VSS nch w=0.175u l=0.06u
MI160 net265 DA net109 VSS nch w=0.175u l=0.06u
MI218-M_u2 QN net098 VSS VSS nch w=0.78u l=0.06u
MI241-M_u2 Q net82 VSS VSS nch w=0.78u l=0.06u
MI243-M_u2 net0124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0122 SA VSS VSS nch w=0.195u l=0.06u
MI214-M_u2 net098 net82 VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 net086 d0 VSS VSS nch w=0.195u l=0.06u
MI29 net82 INCPB net074 VSS nch w=0.15u l=0.06u
MI41 net074 net098 VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SDFXD4 DA DB SA SI SE CP Q QN VDD VSS
MI231 net0147 SE VDD VDD pch w=0.35u l=0.06u
MI250 net82 INCPB net0176 VDD pch w=0.27u l=0.06u
MI251 net0176 net086 VDD VDD pch w=0.27u l=0.06u
MI233 net208 SA net0145 VDD pch w=0.435u l=0.06u
MI232 net0145 DB net0147 VDD pch w=0.255u l=0.06u
MI102 net144 net086 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net144 VDD pch w=0.15u l=0.06u
MI223 net82 INCPB net0171 VDD pch w=0.4u l=0.06u
MI234 net208 net0124 net0148 VDD pch w=0.2u l=0.06u
MI235 net0148 SI VDD VDD pch w=0.2u l=0.06u
MI222 net0171 net086 VDD VDD pch w=0.3u l=0.06u
MI150 net208 DA net162 VDD pch w=0.35u l=0.06u
MI151 net162 net0122 net0147 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net208 VDD pch w=0.35u l=0.06u
MI260-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI256-M_u3 QN net098 VDD VDD pch w=0.52u l=0.06u
MI242-M_u3 QN net098 VDD VDD pch w=0.52u l=0.06u
MI265-M_u3 net0124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0122 SA VDD VDD pch w=0.26u l=0.06u
MI254-M_u3 QN net098 VDD VDD pch w=0.52u l=0.06u
MI255-M_u3 QN net098 VDD VDD pch w=0.52u l=0.06u
MI259-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI258-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI263-M_u3 INCPB CP VDD VDD pch w=0.42u l=0.06u
MI257-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI214-M_u3 net098 net82 VDD VDD pch w=0.46u l=0.06u
MI264-M_u3 INCP INCPB VDD VDD pch w=0.49u l=0.06u
MI123-M_u3 net086 d0 VDD VDD pch w=0.29u l=0.06u
MI38 net82 INCP net070 VDD pch w=0.15u l=0.06u
MI24 net070 net098 VDD VDD pch w=0.15u l=0.06u
MI237 net265 SE net099 VSS nch w=0.15u l=0.06u
MI238 net265 net0122 net096 VSS nch w=0.175u l=0.06u
MI239 net096 DB net093 VSS nch w=0.175u l=0.06u
MI227 net82 INCP net0118 VSS nch w=0.33u l=0.06u
MI248 net82 INCP net0104 VSS nch w=0.245u l=0.06u
MI249 net0104 net086 VSS VSS nch w=0.33u l=0.06u
MI240 net093 net0124 VSS VSS nch w=0.355u l=0.06u
MI119 net79 net086 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net79 VSS nch w=0.15u l=0.06u
MI225 net0118 net086 VSS VSS nch w=0.33u l=0.06u
MI236 net099 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net265 VSS nch w=0.195u l=0.06u
MI163 net109 SA net093 VSS nch w=0.175u l=0.06u
MI160 net265 DA net109 VSS nch w=0.175u l=0.06u
MI260-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI256-M_u2 QN net098 VSS VSS nch w=0.39u l=0.06u
MI242-M_u2 QN net098 VSS VSS nch w=0.39u l=0.06u
MI265-M_u2 net0124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0122 SA VSS VSS nch w=0.195u l=0.06u
MI254-M_u2 QN net098 VSS VSS nch w=0.39u l=0.06u
MI255-M_u2 QN net098 VSS VSS nch w=0.39u l=0.06u
MI259-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI258-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI263-M_u2 INCPB CP VSS VSS nch w=0.31u l=0.06u
MI257-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI214-M_u2 net098 net82 VSS VSS nch w=0.39u l=0.06u
MI264-M_u2 INCP INCPB VSS VSS nch w=0.28u l=0.06u
MI123-M_u2 net086 d0 VSS VSS nch w=0.2u l=0.06u
MI29 net82 INCPB net074 VSS nch w=0.16u l=0.06u
MI41 net074 net098 VSS VSS nch w=0.16u l=0.06u
.ends
.subckt SDFXQD0 DA DB SA SI SE CP Q VDD VSS
MI185 d1 INCPB net278 VDD pch w=0.44u l=0.06u
MI156 net193 SA VDD VDD pch w=0.24u l=0.06u
MI136 net220 Q VDD VDD pch w=0.15u l=0.06u
MI155 net188 net235 VDD VDD pch w=0.24u l=0.06u
MI154 net255 DB net193 VDD pch w=0.24u l=0.06u
MI153 d0 INCP net197 VDD pch w=0.3u l=0.06u
MI152 net197 net233 net199 VDD pch w=0.26u l=0.06u
MI151 net208 SE VDD VDD pch w=0.26u l=0.06u
MI157 net255 DA net188 VDD pch w=0.24u l=0.06u
MI150 net197 net255 net208 VDD pch w=0.26u l=0.06u
MI149 net199 net0110 VDD VDD pch w=0.26u l=0.06u
MI103 d0 INCPB net214 VDD pch w=0.15u l=0.06u
MI186 net278 INCP net220 VDD pch w=0.15u l=0.06u
MI102 net214 d1 VDD VDD pch w=0.15u l=0.06u
MI189-M_u3 net0110 SI VDD VDD pch w=0.15u l=0.06u
MI181-M_u3 Q net278 VDD VDD pch w=0.26u l=0.06u
MI170-M_u3 net235 SA VDD VDD pch w=0.2u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI123-M_u3 d1 d0 VDD VDD pch w=0.34u l=0.06u
MI169-M_u3 net233 SE VDD VDD pch w=0.2u l=0.06u
MI190-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI189-M_u2 net0110 SI VSS VSS nch w=0.15u l=0.06u
MI181-M_u2 Q net278 VSS VSS nch w=0.195u l=0.06u
MI170-M_u2 net235 SA VSS VSS nch w=0.15u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 d1 d0 VSS VSS nch w=0.34u l=0.06u
MI169-M_u2 net233 SE VSS VSS nch w=0.15u l=0.06u
MI190-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI161 net240 SE net264 VSS nch w=0.195u l=0.06u
MI163 net246 net233 VSS VSS nch w=0.195u l=0.06u
MI167 net258 net235 VSS VSS nch w=0.195u l=0.06u
MI164 d0 INCPB net240 VSS nch w=0.2u l=0.06u
MI166 net255 DA net254 VSS nch w=0.195u l=0.06u
MI162 net264 net0110 VSS VSS nch w=0.195u l=0.06u
MI178 d1 INCP net278 VSS nch w=0.22u l=0.06u
MI135 net278 INCPB net267 VSS nch w=0.15u l=0.06u
MI168 net255 DB net258 VSS nch w=0.195u l=0.06u
MI165 net254 SA VSS VSS nch w=0.195u l=0.06u
MI120 d0 INCP net269 VSS nch w=0.15u l=0.06u
MI160 net240 net255 net246 VSS nch w=0.195u l=0.06u
MI119 net269 d1 VSS VSS nch w=0.15u l=0.06u
MI122 net267 Q VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SDFXQD1 DA DB SA SI SE CP Q VDD VSS
MI240 net153 net124 VSS VSS nch w=0.355u l=0.06u
MI119 net145 net146 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net145 VSS nch w=0.15u l=0.06u
MI225 net139 net146 VSS VSS nch w=0.205u l=0.06u
MI237 net160 SE net136 VSS nch w=0.15u l=0.06u
MI236 net136 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net160 VSS nch w=0.195u l=0.06u
MI238 net160 net122 net156 VSS nch w=0.175u l=0.06u
MI163 net126 SA net153 VSS nch w=0.175u l=0.06u
MI160 net160 DA net126 VSS nch w=0.175u l=0.06u
MI239 net156 DB net153 VSS nch w=0.175u l=0.06u
MI227 net94 INCP net139 VSS nch w=0.22u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 net146 d0 VSS VSS nch w=0.195u l=0.06u
MI194-M_u2 net124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net122 SA VSS VSS nch w=0.195u l=0.06u
MI228-M_u2 Q net94 VSS VSS nch w=0.39u l=0.06u
MI193-M_u2 net164 net94 VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI29 net94 INCPB net165 VSS nch w=0.15u l=0.06u
MI41 net165 net164 VSS VSS nch w=0.15u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 net146 d0 VDD VDD pch w=0.26u l=0.06u
MI194-M_u3 net124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net122 SA VDD VDD pch w=0.26u l=0.06u
MI228-M_u3 Q net94 VDD VDD pch w=0.52u l=0.06u
MI193-M_u3 net164 net94 VDD VDD pch w=0.15u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI231 net105 SE VDD VDD pch w=0.35u l=0.06u
MI233 net91 SA net103 VDD pch w=0.435u l=0.06u
MI232 net103 DB net105 VDD pch w=0.255u l=0.06u
MI102 net100 net146 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net100 VDD pch w=0.15u l=0.06u
MI223 net94 INCPB net96 VDD pch w=0.27u l=0.06u
MI234 net91 net124 net88 VDD pch w=0.2u l=0.06u
MI235 net88 SI VDD VDD pch w=0.2u l=0.06u
MI222 net96 net146 VDD VDD pch w=0.27u l=0.06u
MI150 net91 DA net84 VDD pch w=0.35u l=0.06u
MI151 net84 net122 net105 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net91 VDD pch w=0.3u l=0.06u
MI38 net94 INCP net173 VDD pch w=0.15u l=0.06u
MI24 net173 net164 VDD VDD pch w=0.15u l=0.06u
.ends
.subckt SDFXQD2 DA DB SA SI SE CP Q VDD VSS
MI241-M_u3 Q net82 VDD VDD pch w=1.04u l=0.06u
MI243-M_u3 net0124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0122 SA VDD VDD pch w=0.26u l=0.06u
MI214-M_u3 net098 net82 VDD VDD pch w=0.15u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 net086 d0 VDD VDD pch w=0.26u l=0.06u
MI231 net0147 SE VDD VDD pch w=0.35u l=0.06u
MI233 net208 SA net0145 VDD pch w=0.435u l=0.06u
MI232 net0145 DB net0147 VDD pch w=0.255u l=0.06u
MI102 net144 net086 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net144 VDD pch w=0.15u l=0.06u
MI223 net82 INCPB net0171 VDD pch w=0.27u l=0.06u
MI234 net208 net0124 net0148 VDD pch w=0.2u l=0.06u
MI235 net0148 SI VDD VDD pch w=0.2u l=0.06u
MI222 net0171 net086 VDD VDD pch w=0.27u l=0.06u
MI150 net208 DA net162 VDD pch w=0.35u l=0.06u
MI151 net162 net0122 net0147 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net208 VDD pch w=0.3u l=0.06u
MI38 net82 INCP net070 VDD pch w=0.15u l=0.06u
MI24 net070 net098 VDD VDD pch w=0.15u l=0.06u
MI237 net265 SE net099 VSS nch w=0.15u l=0.06u
MI238 net265 net0122 net096 VSS nch w=0.175u l=0.06u
MI239 net096 DB net093 VSS nch w=0.175u l=0.06u
MI227 net82 INCP net0118 VSS nch w=0.22u l=0.06u
MI240 net093 net0124 VSS VSS nch w=0.355u l=0.06u
MI119 net79 net086 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net79 VSS nch w=0.15u l=0.06u
MI225 net0118 net086 VSS VSS nch w=0.205u l=0.06u
MI236 net099 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net265 VSS nch w=0.195u l=0.06u
MI163 net109 SA net093 VSS nch w=0.175u l=0.06u
MI160 net265 DA net109 VSS nch w=0.175u l=0.06u
MI241-M_u2 Q net82 VSS VSS nch w=0.78u l=0.06u
MI243-M_u2 net0124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0122 SA VSS VSS nch w=0.195u l=0.06u
MI214-M_u2 net098 net82 VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 net086 d0 VSS VSS nch w=0.195u l=0.06u
MI29 net82 INCPB net074 VSS nch w=0.15u l=0.06u
MI41 net074 net098 VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SDFXQD4 DA DB SA SI SE CP Q VDD VSS
MI231 net0147 SE VDD VDD pch w=0.35u l=0.06u
MI250 net82 INCPB net0176 VDD pch w=0.27u l=0.06u
MI251 net0176 net086 VDD VDD pch w=0.27u l=0.06u
MI233 net208 SA net0145 VDD pch w=0.435u l=0.06u
MI232 net0145 DB net0147 VDD pch w=0.255u l=0.06u
MI102 net144 net086 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net144 VDD pch w=0.15u l=0.06u
MI223 net82 INCPB net0171 VDD pch w=0.4u l=0.06u
MI234 net208 net0124 net0148 VDD pch w=0.2u l=0.06u
MI235 net0148 SI VDD VDD pch w=0.2u l=0.06u
MI222 net0171 net086 VDD VDD pch w=0.3u l=0.06u
MI150 net208 DA net162 VDD pch w=0.35u l=0.06u
MI151 net162 net0122 net0147 VDD pch w=0.35u l=0.06u
MI153 d0 INCP net208 VDD pch w=0.35u l=0.06u
MI260-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI264-M_u3 INCP INCPB VDD VDD pch w=0.49u l=0.06u
MI263-M_u3 INCPB CP VDD VDD pch w=0.42u l=0.06u
MI265-M_u3 net0124 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0122 SA VDD VDD pch w=0.26u l=0.06u
MI259-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI258-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI257-M_u3 Q net82 VDD VDD pch w=0.52u l=0.06u
MI214-M_u3 net098 net82 VDD VDD pch w=0.15u l=0.06u
MI123-M_u3 net086 d0 VDD VDD pch w=0.29u l=0.06u
MI38 net82 INCP net070 VDD pch w=0.15u l=0.06u
MI24 net070 net098 VDD VDD pch w=0.15u l=0.06u
MI237 net265 SE net099 VSS nch w=0.15u l=0.06u
MI238 net265 net0122 net096 VSS nch w=0.175u l=0.06u
MI239 net096 DB net093 VSS nch w=0.175u l=0.06u
MI227 net82 INCP net0118 VSS nch w=0.33u l=0.06u
MI248 net82 INCP net0104 VSS nch w=0.245u l=0.06u
MI249 net0104 net086 VSS VSS nch w=0.33u l=0.06u
MI240 net093 net0124 VSS VSS nch w=0.355u l=0.06u
MI119 net79 net086 VSS VSS nch w=0.15u l=0.06u
MI120 d0 INCP net79 VSS nch w=0.15u l=0.06u
MI225 net0118 net086 VSS VSS nch w=0.33u l=0.06u
MI236 net099 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net265 VSS nch w=0.195u l=0.06u
MI163 net109 SA net093 VSS nch w=0.175u l=0.06u
MI160 net265 DA net109 VSS nch w=0.175u l=0.06u
MI260-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI264-M_u2 INCP INCPB VSS VSS nch w=0.28u l=0.06u
MI263-M_u2 INCPB CP VSS VSS nch w=0.31u l=0.06u
MI265-M_u2 net0124 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0122 SA VSS VSS nch w=0.195u l=0.06u
MI259-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI258-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI257-M_u2 Q net82 VSS VSS nch w=0.39u l=0.06u
MI214-M_u2 net098 net82 VSS VSS nch w=0.16u l=0.06u
MI123-M_u2 net086 d0 VSS VSS nch w=0.2u l=0.06u
MI29 net82 INCPB net074 VSS nch w=0.16u l=0.06u
MI41 net074 net098 VSS VSS nch w=0.16u l=0.06u
.ends
.subckt SEDFCND0 E SE CP SI D CDN Q QN VDD VSS
MI191-M_u2 net78 CDN VDD VDD pch w=0.4u l=0.06u
MI191-M_u1 net78 net139 VDD VDD pch w=0.4u l=0.06u
MI178 net156 net134 net139 VDD pch w=0.15u l=0.06u
MI153 d0 net134 net87 VDD pch w=0.25u l=0.06u
MI150 net87 D net96 VDD pch w=0.47u l=0.06u
MI233 net87 E net90 VDD pch w=0.375u l=0.06u
MI151 net96 net130 net92 VDD pch w=0.32u l=0.06u
MI179 d1 INCPB net139 VDD pch w=0.39u l=0.06u
MI232 net90 net156 net92 VDD pch w=0.255u l=0.06u
MI234 net87 net120 net89 VDD pch w=0.15u l=0.06u
MI231 net92 SE VDD VDD pch w=0.32u l=0.06u
MI235 net89 SI VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net119 VDD pch w=0.15u l=0.06u
MI102 net119 d1 VDD VDD pch w=0.15u l=0.06u
MI101 net119 CDN VDD VDD pch w=0.15u l=0.06u
MI192-M_u3 net130 E VDD VDD pch w=0.2u l=0.06u
MI189-M_u3 QN net156 VDD VDD pch w=0.26u l=0.06u
MI177-M_u3 net156 net78 VDD VDD pch w=0.2u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI188-M_u3 Q net78 VDD VDD pch w=0.26u l=0.06u
MI230-M_u3 net120 SE VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 net134 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI191-M_u4 XI191-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI191-M_u3 net78 net139 XI191-net6 VSS nch w=0.23u l=0.06u
MI192-M_u2 net130 E VSS VSS nch w=0.15u l=0.06u
MI189-M_u2 QN net156 VSS VSS nch w=0.195u l=0.06u
MI177-M_u2 net156 net78 VSS VSS nch w=0.15u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI188-M_u2 Q net78 VSS VSS nch w=0.195u l=0.06u
MI230-M_u2 net120 SE VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 net134 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI173 net156 INCPB net139 VSS nch w=0.15u l=0.06u
MI119 net167 d1 net166 VSS nch w=0.15u l=0.06u
MI240 net154 net120 VSS VSS nch w=0.355u l=0.06u
MI120 d0 net134 net167 VSS nch w=0.15u l=0.06u
MI236 net151 SI VSS VSS nch w=0.15u l=0.06u
MI239 net145 net156 net154 VSS nch w=0.175u l=0.06u
MI237 net152 SE net151 VSS nch w=0.15u l=0.06u
MI163 net149 E net154 VSS nch w=0.355u l=0.06u
MI238 net152 net130 net145 VSS nch w=0.175u l=0.06u
MI160 net152 D net149 VSS nch w=0.26u l=0.06u
MI174 d1 net134 net139 VSS nch w=0.17u l=0.06u
MI164 d0 INCPB net152 VSS nch w=0.34u l=0.06u
MI118 net166 CDN VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFCND1 E SE CP SI D CDN Q QN VDD VSS
MI237 net076 SE net0102 VSS nch w=0.15u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI188-M_u2 Q net077 VSS VSS nch w=0.39u l=0.06u
MI189-M_u2 QN net0124 VSS VSS nch w=0.39u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.195u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI193-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MI192-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 net0122 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI191-M_u4 XI191-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI191-M_u3 net077 net76 XI191-net6 VSS nch w=0.23u l=0.06u
MI188-M_u3 Q net077 VDD VDD pch w=0.52u l=0.06u
MI189-M_u3 QN net0124 VDD VDD pch w=0.52u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI193-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MI192-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 net0122 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.25u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.15u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.15u l=0.06u
MI191-M_u2 net077 CDN VDD VDD pch w=0.4u l=0.06u
MI191-M_u1 net077 net76 VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SEDFCND2 E SE CP SI D CDN Q QN VDD VSS
MI237 net076 SE net0102 VSS nch w=0.15u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI193-M_u2 QN net0124 VSS VSS nch w=0.39u l=0.06u
MI197-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MI194-M_u2 Q net077 VSS VSS nch w=0.39u l=0.06u
MI195-M_u2 Q net077 VSS VSS nch w=0.39u l=0.06u
MI192-M_u2 QN net0124 VSS VSS nch w=0.39u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.195u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI198-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 net0122 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI196-M_u4 XI196-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI196-M_u3 net077 net76 XI196-net6 VSS nch w=0.23u l=0.06u
MI193-M_u3 QN net0124 VDD VDD pch w=0.52u l=0.06u
MI197-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MI194-M_u3 Q net077 VDD VDD pch w=0.52u l=0.06u
MI195-M_u3 Q net077 VDD VDD pch w=0.52u l=0.06u
MI192-M_u3 QN net0124 VDD VDD pch w=0.52u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI198-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 net0122 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.25u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.15u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.15u l=0.06u
MI196-M_u2 net077 CDN VDD VDD pch w=0.4u l=0.06u
MI196-M_u1 net077 net76 VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SEDFCND4 E SE CP SI D CDN Q QN VDD VSS
MI237 net076 SE net0102 VSS nch w=0.15u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI188-M_u2 Q net077 VSS VSS nch w=1.56u l=0.06u
MI189-M_u2 QN net0124 VSS VSS nch w=1.56u l=0.06u
MI201-M_u2 net0122 INCPB VSS VSS nch w=0.39u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.19u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI203-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MI202-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI183-M_u4 XI183-net6 net76 VSS VSS nch w=0.225u l=0.06u
MI183-M_u3 net077 CDN XI183-net6 VSS nch w=0.225u l=0.06u
MI197-M_u4 XI197-net6 net76 VSS VSS nch w=0.225u l=0.06u
MI197-M_u3 net077 CDN XI197-net6 VSS nch w=0.225u l=0.06u
MI188-M_u3 Q net077 VDD VDD pch w=2.08u l=0.06u
MI189-M_u3 QN net0124 VDD VDD pch w=2.08u l=0.06u
MI201-M_u3 net0122 INCPB VDD VDD pch w=0.52u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI203-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MI202-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.34u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.15u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.15u l=0.06u
MI183-M_u2 net077 net76 VDD VDD pch w=0.52u l=0.06u
MI183-M_u1 net077 CDN VDD VDD pch w=0.52u l=0.06u
MI197-M_u2 net077 net76 VDD VDD pch w=0.52u l=0.06u
MI197-M_u1 net077 CDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SEDFCNQD0 E SE CP SI D CDN Q VDD VSS
MI191-M_u2 net76 CDN VDD VDD pch w=0.4u l=0.06u
MI191-M_u1 net76 net156 VDD VDD pch w=0.4u l=0.06u
MI178 net149 net124 net156 VDD pch w=0.15u l=0.06u
MI179 d1 INCPB net156 VDD pch w=0.39u l=0.06u
MI153 d0 net124 net85 VDD pch w=0.25u l=0.06u
MI150 net85 D net91 VDD pch w=0.47u l=0.06u
MI233 net85 E net88 VDD pch w=0.2u l=0.06u
MI151 net91 net120 net90 VDD pch w=0.32u l=0.06u
MI103 d0 INCPB net117 VDD pch w=0.15u l=0.06u
MI232 net88 net149 net90 VDD pch w=0.2u l=0.06u
MI234 net85 net118 net87 VDD pch w=0.15u l=0.06u
MI231 net90 SE VDD VDD pch w=0.32u l=0.06u
MI235 net87 SI VDD VDD pch w=0.15u l=0.06u
MI102 net117 d1 VDD VDD pch w=0.15u l=0.06u
MI101 net117 CDN VDD VDD pch w=0.15u l=0.06u
MI188-M_u3 Q net76 VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 net124 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI197-M_u3 net120 E VDD VDD pch w=0.2u l=0.06u
MI198-M_u3 net118 SE VDD VDD pch w=0.2u l=0.06u
MI177-M_u3 net149 net76 VDD VDD pch w=0.2u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI191-M_u4 XI191-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI191-M_u3 net76 net156 XI191-net6 VSS nch w=0.23u l=0.06u
MI188-M_u2 Q net76 VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 net124 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI197-M_u2 net120 E VSS VSS nch w=0.15u l=0.06u
MI198-M_u2 net118 SE VSS VSS nch w=0.15u l=0.06u
MI177-M_u2 net149 net76 VSS VSS nch w=0.15u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI173 net149 INCPB net156 VSS nch w=0.15u l=0.06u
MI119 net163 d1 net169 VSS nch w=0.15u l=0.06u
MI120 d0 net124 net163 VSS nch w=0.15u l=0.06u
MI174 d1 net124 net156 VSS nch w=0.17u l=0.06u
MI240 net147 net118 VSS VSS nch w=0.355u l=0.06u
MI236 net151 SI VSS VSS nch w=0.15u l=0.06u
MI239 net148 net149 net147 VSS nch w=0.175u l=0.06u
MI237 net145 SE net151 VSS nch w=0.15u l=0.06u
MI163 net135 E net147 VSS nch w=0.355u l=0.06u
MI238 net145 net120 net148 VSS nch w=0.175u l=0.06u
MI160 net145 D net135 VSS nch w=0.26u l=0.06u
MI164 d0 INCPB net145 VSS nch w=0.34u l=0.06u
MI118 net169 CDN VSS VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFCNQD1 E SE CP SI D CDN Q VDD VSS
MI237 net076 SE net0102 VSS nch w=0.15u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI188-M_u2 Q net077 VSS VSS nch w=0.39u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.195u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI193-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MI192-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 net0122 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI191-M_u4 XI191-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI191-M_u3 net077 net76 XI191-net6 VSS nch w=0.23u l=0.06u
MI188-M_u3 Q net077 VDD VDD pch w=0.52u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI193-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MI192-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 net0122 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.25u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.2u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.2u l=0.06u
MI191-M_u2 net077 CDN VDD VDD pch w=0.4u l=0.06u
MI191-M_u1 net077 net76 VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SEDFCNQD2 E SE CP SI D CDN Q VDD VSS
MI237 net076 SE net0102 VSS nch w=0.19u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.19u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI188-M_u2 Q net077 VSS VSS nch w=0.78u l=0.06u
MI193-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.195u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI194-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 net0122 INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI192-M_u4 XI192-net6 CDN VSS VSS nch w=0.23u l=0.06u
MI192-M_u3 net077 net76 XI192-net6 VSS nch w=0.23u l=0.06u
MI188-M_u3 Q net077 VDD VDD pch w=1.04u l=0.06u
MI193-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI194-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 net0122 INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.25u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.26u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.26u l=0.06u
MI192-M_u2 net077 CDN VDD VDD pch w=0.4u l=0.06u
MI192-M_u1 net077 net76 VDD VDD pch w=0.4u l=0.06u
.ends
.subckt SEDFCNQD4 E SE CP SI D CDN Q VDD VSS
MI237 net076 SE net0102 VSS nch w=0.15u l=0.06u
MI174 d1 net0122 net76 VSS nch w=0.17u l=0.06u
MI173 net0124 INCPB net76 VSS nch w=0.15u l=0.06u
MI118 net92 CDN VSS VSS nch w=0.15u l=0.06u
MI119 net95 d1 net92 VSS nch w=0.15u l=0.06u
MI120 d0 net0122 net95 VSS nch w=0.15u l=0.06u
MI240 net096 net0126 VSS VSS nch w=0.355u l=0.06u
MI236 net0102 SI VSS VSS nch w=0.15u l=0.06u
MI164 d0 INCPB net076 VSS nch w=0.34u l=0.06u
MI163 net085 E net096 VSS nch w=0.355u l=0.06u
MI160 net076 D net085 VSS nch w=0.26u l=0.06u
MI238 net076 net0103 net099 VSS nch w=0.175u l=0.06u
MI239 net099 net0124 net096 VSS nch w=0.175u l=0.06u
MI188-M_u2 Q net077 VSS VSS nch w=1.56u l=0.06u
MI196-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI198-M_u2 net0103 E VSS VSS nch w=0.195u l=0.06u
MI177-M_u2 net0124 net077 VSS VSS nch w=0.19u l=0.06u
MI190-M_u2 d1 d0 VSS VSS nch w=0.21u l=0.06u
MI230-M_u2 net0126 SE VSS VSS nch w=0.195u l=0.06u
MI197-M_u2 net0122 INCPB VSS VSS nch w=0.39u l=0.06u
MI183-M_u4 XI183-net6 net76 VSS VSS nch w=0.23u l=0.06u
MI183-M_u3 net077 CDN XI183-net6 VSS nch w=0.23u l=0.06u
MI194-M_u4 XI194-net6 net76 VSS VSS nch w=0.23u l=0.06u
MI194-M_u3 net077 CDN XI194-net6 VSS nch w=0.23u l=0.06u
MI188-M_u3 Q net077 VDD VDD pch w=2.08u l=0.06u
MI196-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI198-M_u3 net0103 E VDD VDD pch w=0.26u l=0.06u
MI177-M_u3 net0124 net077 VDD VDD pch w=0.26u l=0.06u
MI190-M_u3 d1 d0 VDD VDD pch w=0.21u l=0.06u
MI230-M_u3 net0126 SE VDD VDD pch w=0.26u l=0.06u
MI197-M_u3 net0122 INCPB VDD VDD pch w=0.52u l=0.06u
MI231 net0153 SE VDD VDD pch w=0.32u l=0.06u
MI233 net0148 E net0151 VDD pch w=0.375u l=0.06u
MI101 net83 CDN VDD VDD pch w=0.15u l=0.06u
MI178 net0124 net0122 net76 VDD pch w=0.15u l=0.06u
MI102 net83 d1 VDD VDD pch w=0.15u l=0.06u
MI103 d0 INCPB net83 VDD pch w=0.15u l=0.06u
MI150 net0148 D net0144 VDD pch w=0.47u l=0.06u
MI179 d1 INCPB net76 VDD pch w=0.39u l=0.06u
MI232 net0151 net0124 net0153 VDD pch w=0.255u l=0.06u
MI151 net0144 net0103 net0153 VDD pch w=0.32u l=0.06u
MI153 d0 net0122 net0148 VDD pch w=0.34u l=0.06u
MI234 net0148 net0126 net0145 VDD pch w=0.2u l=0.06u
MI235 net0145 SI VDD VDD pch w=0.2u l=0.06u
MI183-M_u2 net077 net76 VDD VDD pch w=0.52u l=0.06u
MI183-M_u1 net077 CDN VDD VDD pch w=0.52u l=0.06u
MI194-M_u2 net077 net76 VDD VDD pch w=0.52u l=0.06u
MI194-M_u1 net077 CDN VDD VDD pch w=0.52u l=0.06u
.ends
.subckt SEDFD0 E SE CP SI D Q QN VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.26u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI228-M_u3 QN SLO VDD VDD pch w=0.26u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.2u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.195u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI228-M_u2 QN SLO VSS VSS nch w=0.195u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.15u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFD1 E SE CP SI D Q QN VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFD2 E SE CP SI D Q QN VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI236-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI237-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI236-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI237-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFD4 E SE CP SI D Q QN VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI236-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI237-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI238-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI239-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI243-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI240-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI241-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI245-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI242-M_u3 SLO SLI VDD VDD pch w=0.52u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MI244-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI236-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI237-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI238-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI239-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI243-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI240-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI241-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI245-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI242-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MI244-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFKCND0 SI D E SE CP CN Q QN VDD VSS
MI146 net84 CN VSS VSS nch w=0.15u l=0.06u
MI144 net189 D net086 VSS nch w=0.37u l=0.06u
MI145 net086 E net84 VSS nch w=0.15u l=0.06u
MI143 net95 net185 net84 VSS nch w=0.37u l=0.06u
MI113 net189 net101 net95 VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI64 net102 net93 VSS VSS nch w=0.275u l=0.06u
MI65 net193 net163 net102 VSS nch w=0.275u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI135-M_u2 Q net156 VSS VSS nch w=0.195u l=0.06u
MI148-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI48-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.15u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI138-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI149-M_u2 net185 net156 VSS VSS nch w=0.15u l=0.06u
MI130-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI147-M_u2 QN net185 VSS VSS nch w=0.195u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.15u l=0.06u
MI135-M_u3 Q net156 VDD VDD pch w=0.26u l=0.06u
MI148-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI48-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.2u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI138-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI149-M_u3 net185 net156 VDD VDD pch w=0.2u l=0.06u
MI130-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI147-M_u3 QN net185 VDD VDD pch w=0.26u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.2u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI140 net0150 net185 VDD VDD pch w=0.21u l=0.06u
MI142 net189 CN VDD VDD pch w=0.2u l=0.06u
MI141 net189 E net0150 VDD pch w=0.21u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI50 net174 SE VDD VDD pch w=0.355u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.15u l=0.06u
MI51 net145 net163 net174 VDD pch w=0.175u l=0.06u
MI52 net72 SI VDD VDD pch w=0.15u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
MI139 net189 D net151 VDD pch w=0.34u l=0.06u
.ends
.subckt SEDFKCND1 SI D E SE CP CN Q QN VDD VSS
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI153 net189 net101 net087 VSS nch w=0.37u l=0.06u
MI154 net087 net185 net84 VSS nch w=0.37u l=0.06u
MI112 net84 CN VSS VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI152 net87 E net84 VSS nch w=0.19u l=0.06u
MI143-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI157-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI158-M_u2 net185 net156 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI132-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI143-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI157-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI158-M_u3 net185 net156 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI132-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI149 net0151 net185 VDD VDD pch w=0.21u l=0.06u
MI150 net189 E net0151 VDD pch w=0.21u l=0.06u
MI146 net189 D net151 VDD pch w=0.34u l=0.06u
MI155 net189 CN VDD VDD pch w=0.36u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.15u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.15u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
.ends
.subckt SEDFKCND2 SI D E SE CP CN Q QN VDD VSS
MI158 net84 CN VSS VSS nch w=0.37u l=0.06u
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI153 net189 net101 net087 VSS nch w=0.37u l=0.06u
MI154 net087 net185 net84 VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI152 net87 E net84 VSS nch w=0.19u l=0.06u
MI156-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI157-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI162-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI160-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI161-M_u2 net185 net156 VSS VSS nch w=0.195u l=0.06u
MI130-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI132-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI156-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI157-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI162-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI160-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI161-M_u3 net185 net156 VDD VDD pch w=0.26u l=0.06u
MI130-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI132-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI149 net0151 net185 VDD VDD pch w=0.21u l=0.06u
MI150 net189 E net0151 VDD pch w=0.21u l=0.06u
MI146 net189 D net151 VDD pch w=0.34u l=0.06u
MI155 net189 CN VDD VDD pch w=0.36u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.175u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.175u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
.ends
.subckt SEDFKCND4 SI D E SE CP CN Q QN VDD VSS
MI158 net84 CN VSS VSS nch w=0.37u l=0.06u
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI153 net189 net101 net087 VSS nch w=0.37u l=0.06u
MI154 net087 net185 net84 VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI152 net87 E net84 VSS nch w=0.19u l=0.06u
MI156-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI159-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI157-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI160-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI161-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI162-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI163-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI169-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI166-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI164-M_u2 net185 net156 VSS VSS nch w=0.78u l=0.06u
MI130-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI132-M_u2 QN net185 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI156-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI159-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI157-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI160-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI161-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI162-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI163-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI169-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI166-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI164-M_u3 net185 net156 VDD VDD pch w=1.04u l=0.06u
MI130-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI132-M_u3 QN net185 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI149 net0151 net185 VDD VDD pch w=0.21u l=0.06u
MI150 net189 E net0151 VDD pch w=0.21u l=0.06u
MI146 net189 D net151 VDD pch w=0.34u l=0.06u
MI155 net189 CN VDD VDD pch w=0.36u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.41u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.175u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.175u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
.ends
.subckt SEDFKCNQD0 SI D E SE CP CN Q VDD VSS
MI145-M_u2 net081 SI VSS VSS nch w=0.15u l=0.06u
MI148-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI146-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.34u l=0.06u
MI130-M_u2 Q net83 VSS VSS nch w=0.375u l=0.06u
MI147-M_u2 net101 E VSS VSS nch w=0.15u l=0.06u
MI141 net95 Q net84 VSS nch w=0.195u l=0.06u
MI143 net099 E net84 VSS nch w=0.17u l=0.06u
MI144 net84 CN VSS VSS nch w=0.15u l=0.06u
MI142 net189 D net099 VSS nch w=0.195u l=0.06u
MI113 net189 net101 net95 VSS nch w=0.195u l=0.06u
MI29 net83 INCPB net083 VSS nch w=0.15u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.18u l=0.06u
MI39 net083 Q VSS VSS nch w=0.15u l=0.06u
MI64 net102 net93 VSS VSS nch w=0.195u l=0.06u
MI65 net193 net189 net102 VSS nch w=0.195u l=0.06u
MI62 net193 SE net129 VSS nch w=0.195u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.23u l=0.06u
MI63 net129 net081 VSS VSS nch w=0.195u l=0.06u
MI145-M_u3 net081 SI VDD VDD pch w=0.2u l=0.06u
MI148-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.29u l=0.06u
MI146-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.34u l=0.06u
MI130-M_u3 Q net83 VDD VDD pch w=0.52u l=0.06u
MI147-M_u3 net101 E VDD VDD pch w=0.2u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.26u l=0.06u
MI139 net189 E net0146 VDD pch w=0.17u l=0.06u
MI138 net0146 Q VDD VDD pch w=0.17u l=0.06u
MI137 net189 D net151 VDD pch w=0.26u l=0.06u
MI38 net83 INCP net091 VDD pch w=0.15u l=0.06u
MI24 net091 Q VDD VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.43u l=0.06u
MI50 net174 SE VDD VDD pch w=0.255u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.3u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.255u l=0.06u
MI51 net145 net189 net174 VDD pch w=0.255u l=0.06u
MI52 net72 net081 VDD VDD pch w=0.255u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
MI140 net189 CN VDD VDD pch w=0.2u l=0.06u
.ends
.subckt SEDFKCNQD1 SI D E SE CP CN Q VDD VSS
MI149 net95 net185 net84 VSS nch w=0.37u l=0.06u
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI151 net84 CN VSS VSS nch w=0.37u l=0.06u
MI150 net87 E net84 VSS nch w=0.19u l=0.06u
MI113 net189 net101 net95 VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI143-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI152-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI153-M_u2 net185 net156 VSS VSS nch w=0.15u l=0.06u
MI130-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI143-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI152-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI153-M_u3 net185 net156 VDD VDD pch w=0.15u l=0.06u
MI130-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI147 net189 E net0150 VDD pch w=0.21u l=0.06u
MI146 net0150 net185 VDD VDD pch w=0.21u l=0.06u
MI145 net189 D net151 VDD pch w=0.34u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.26u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.175u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.175u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
MI148 net189 CN VDD VDD pch w=0.36u l=0.06u
.ends
.subckt SEDFKCNQD2 SI D E SE CP CN Q VDD VSS
MI146 net088 net185 net84 VSS nch w=0.37u l=0.06u
MI147 net87 E net84 VSS nch w=0.19u l=0.06u
MI145 net189 net101 net088 VSS nch w=0.37u l=0.06u
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI154 net84 CN VSS VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI135-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI143-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI155-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI156-M_u2 net185 net156 VSS VSS nch w=0.15u l=0.06u
MI152-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI135-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI143-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI155-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI156-M_u3 net185 net156 VDD VDD pch w=0.15u l=0.06u
MI152-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI150 net189 E net0151 VDD pch w=0.21u l=0.06u
MI149 net0151 net185 VDD VDD pch w=0.21u l=0.06u
MI148 net189 D net151 VDD pch w=0.34u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.175u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.175u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
MI151 net189 CN VDD VDD pch w=0.36u l=0.06u
.ends
.subckt SEDFKCNQD4 SI D E SE CP CN Q VDD VSS
MI146 net088 net185 net84 VSS nch w=0.37u l=0.06u
MI147 net87 E net84 VSS nch w=0.19u l=0.06u
MI145 net189 net101 net088 VSS nch w=0.37u l=0.06u
MI114 net189 D net87 VSS nch w=0.37u l=0.06u
MI154 net84 CN VSS VSS nch w=0.37u l=0.06u
MI127 net176 INCP net83 VSS nch w=0.21u l=0.06u
MI128 net185 INCPB net83 VSS nch w=0.15u l=0.06u
MI141 net193 net93 net92 VSS nch w=0.21u l=0.06u
MI65 net92 net163 VSS VSS nch w=0.39u l=0.06u
MI62 net193 SE net129 VSS nch w=0.15u l=0.06u
MI101 net175 INCP net123 VSS nch w=0.15u l=0.06u
MI102 net123 net176 VSS VSS nch w=0.15u l=0.06u
MI83 net175 INCPB net193 VSS nch w=0.25u l=0.06u
MI63 net129 SI VSS VSS nch w=0.15u l=0.06u
MI135-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI155-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI158-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI153-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI157-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI156-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI161-M_u2 net185 net156 VSS VSS nch w=0.15u l=0.06u
MI45-M_u2 net93 SE VSS VSS nch w=0.195u l=0.06u
MI42-M_u2 net176 net175 VSS VSS nch w=0.21u l=0.06u
MI105-M_u2 net163 net189 VSS VSS nch w=0.22u l=0.06u
MI152-M_u2 net156 net83 VSS VSS nch w=0.39u l=0.06u
MI131-M_u2 Q net156 VSS VSS nch w=0.39u l=0.06u
MI106-M_u2 net101 E VSS VSS nch w=0.195u l=0.06u
MI135-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI155-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI158-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI153-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI157-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI156-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI161-M_u3 net185 net156 VDD VDD pch w=0.15u l=0.06u
MI45-M_u3 net93 SE VDD VDD pch w=0.255u l=0.06u
MI42-M_u3 net176 net175 VDD VDD pch w=0.23u l=0.06u
MI105-M_u3 net163 net189 VDD VDD pch w=0.52u l=0.06u
MI152-M_u3 net156 net83 VDD VDD pch w=0.52u l=0.06u
MI131-M_u3 Q net156 VDD VDD pch w=0.52u l=0.06u
MI106-M_u3 net101 E VDD VDD pch w=0.26u l=0.06u
MI142 net145 SE net92 VDD pch w=0.355u l=0.06u
MI108 net151 net101 VDD VDD pch w=0.34u l=0.06u
MI150 net189 E net0151 VDD pch w=0.21u l=0.06u
MI149 net0151 net185 VDD VDD pch w=0.21u l=0.06u
MI148 net189 D net151 VDD pch w=0.34u l=0.06u
MI133 net185 INCP net83 VDD pch w=0.15u l=0.06u
MI134 net176 INCPB net83 VDD pch w=0.33u l=0.06u
MI82 net175 INCP net145 VDD pch w=0.34u l=0.06u
MI53 net145 net93 net72 VDD pch w=0.175u l=0.06u
MI51 net92 net163 VDD VDD pch w=0.52u l=0.06u
MI52 net72 SI VDD VDD pch w=0.175u l=0.06u
MI99 net175 INCPB net190 VDD pch w=0.15u l=0.06u
MI100 net190 net176 VDD VDD pch w=0.15u l=0.06u
MI151 net189 CN VDD VDD pch w=0.36u l=0.06u
.ends
.subckt SEDFQD0 E SE CP SI D Q VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.26u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.2u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.195u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.15u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQD1 E SE CP SI D Q VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQD2 E SE CP SI D Q VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI236-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI236-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQD4 E SE CP SI D Q VDD VSS
MI218-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI242-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI244-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI236-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI238-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI239-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MI243-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI218-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI242-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI244-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI236-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI238-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI239-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MI243-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQND0 E SE CP SI D QN VDD VSS
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI228-M_u3 QN SLO VDD VDD pch w=0.26u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.2u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI228-M_u2 QN SLO VSS VSS nch w=0.195u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.15u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQND1 E SE CP SI D QN VDD VSS
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQND2 E SE CP SI D QN VDD VSS
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI237-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI225-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MU84-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI237-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI225-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MU84-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQND4 E SE CP SI D QN VDD VSS
MI243-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI245-M_u3 SLO SLI VDD VDD pch w=0.52u l=0.06u
MI224-M_u3 net0123 SI VDD VDD pch w=0.15u l=0.06u
MI237-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI240-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI241-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI242-M_u3 SLO SLI VDD VDD pch w=0.52u l=0.06u
MI235-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI170-M_u3 net316 E VDD VDD pch w=0.26u l=0.06u
MI169-M_u3 net318 SE VDD VDD pch w=0.26u l=0.06u
MI244-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI231 net094 SLO VDD VDD pch w=0.2u l=0.06u
MI232 SLI INCP net094 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.38u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI149 net167 net0123 VDD VDD pch w=0.2u l=0.06u
MI150 net208 net314 net162 VDD pch w=0.26u l=0.06u
MI157 net314 D net161 VDD pch w=0.26u l=0.06u
MI151 net162 SE VDD VDD pch w=0.26u l=0.06u
MI152 net208 net318 net167 VDD pch w=0.2u l=0.06u
MI153 MLI INCP net208 VDD pch w=0.36u l=0.06u
MI154 net314 E net173 VDD pch w=0.26u l=0.06u
MI155 net161 net316 VDD VDD pch w=0.26u l=0.06u
MI156 net173 SLO VDD VDD pch w=0.26u l=0.06u
MI243-M_u2 INCPB CP VSS VSS nch w=0.39u l=0.06u
MI245-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI224-M_u2 net0123 SI VSS VSS nch w=0.15u l=0.06u
MI237-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI240-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI241-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI242-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI235-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI170-M_u2 net316 E VSS VSS nch w=0.195u l=0.06u
MI169-M_u2 net318 SE VSS VSS nch w=0.18u l=0.06u
MI244-M_u2 INCP INCPB VSS VSS nch w=0.39u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI233 net0135 SLO VSS VSS nch w=0.15u l=0.06u
MI234 SLI INCPB net0135 VSS nch w=0.15u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI162 net112 net0123 VSS VSS nch w=0.15u l=0.06u
MI168 net314 net316 net95 VSS nch w=0.195u l=0.06u
MI167 net95 SLO VSS VSS nch w=0.195u l=0.06u
MI166 net314 D net101 VSS nch w=0.195u l=0.06u
MI165 net101 E VSS VSS nch w=0.195u l=0.06u
MI164 MLI INCPB net265 VSS nch w=0.15u l=0.06u
MI163 net109 net318 VSS VSS nch w=0.16u l=0.06u
MI160 net265 net314 net109 VSS nch w=0.16u l=0.06u
MI161 net265 SE net112 VSS nch w=0.15u l=0.06u
.ends
.subckt SEDFQNXD0 E SE CP SI D QN VDD VSS
MI79 net110 E net107 VSS nch w=0.15u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI255 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.15u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.15u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 QN SLO VSS VSS nch w=0.195u l=0.06u
MI257-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI256 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.2u l=0.06u
MI77 VDD E net110 VDD pch w=0.2u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.2u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 QN SLO VDD VDD pch w=0.26u l=0.06u
MI257-M_u3 d5 SLO VDD VDD pch w=0.2u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.19u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQNXD1 E SE CP SI D QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI255 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI257-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI256 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI257-M_u3 d5 SLO VDD VDD pch w=0.2u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.19u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQNXD2 E SE CP SI D QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI255 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI258-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI212-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI257-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI256 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI258-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI212-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI257-M_u3 d5 SLO VDD VDD pch w=0.15u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQNXD4 E SE CP SI D QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI255 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI258-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI259-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI260-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI262-M_u2 INCPB CP VSS VSS nch w=0.29u l=0.06u
MI212-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI257-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI264-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI261-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI265-M_u2 INCP INCPB VSS VSS nch w=0.29u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI256 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI258-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI259-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI260-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI262-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI212-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI257-M_u3 d5 SLO VDD VDD pch w=0.2u l=0.06u
MI264-M_u3 SLO SLI VDD VDD pch w=0.52u l=0.06u
MI261-M_u3 SLO SLI VDD VDD pch w=0.52u l=0.06u
MI265-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQXD0 E SE CP SI D Q VDD VSS
MI79 net110 E net107 VSS nch w=0.15u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI244 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.15u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.15u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI249-M_u2 Q SLI VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI256-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI243 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.2u l=0.06u
MI77 VDD E net110 VDD pch w=0.2u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.2u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI249-M_u3 Q SLI VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI256-M_u3 d5 SLO VDD VDD pch w=0.15u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQXD1 E SE CP SI D Q VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI244 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI256-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI243 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI256-M_u3 d5 SLO VDD VDD pch w=0.15u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQXD2 E SE CP SI D Q VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI244 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI255-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI256-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI243 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI255-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI256-M_u3 d5 SLO VDD VDD pch w=0.15u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFQXD4 E SE CP SI D Q VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 d5 net108 net104 VSS nch w=0.195u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI244 SLI INCPB d5 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI255-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI268-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI265-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI259-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI260-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI271-M_u2 INCPB CP VSS VSS nch w=0.29u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI270-M_u2 INCP INCPB VSS VSS nch w=0.29u l=0.06u
MI267-M_u2 d5 SLO VSS VSS nch w=0.15u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 d5 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI243 SLI INCP d5 VDD pch w=0.15u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI255-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI268-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI265-M_u3 SLO SLI VDD VDD pch w=0.15u l=0.06u
MI259-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI260-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI271-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI270-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI267-M_u3 d5 SLO VDD VDD pch w=0.15u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFXD0 E SE CP SI D Q QN VDD VSS
MI79 net110 E net107 VSS nch w=0.15u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 net0109 net108 net104 VSS nch w=0.195u l=0.06u
MI251 SLI INCPB net096 VSS nch w=0.15u l=0.06u
MI250 net096 SLO VSS VSS nch w=0.15u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.15u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.15u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.195u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.15u l=0.06u
MI256-M_u2 QN SLO VSS VSS nch w=0.15u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MI257-M_u2 net0109 SLO VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 net0109 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI253 net0143 SLO VDD VDD pch w=0.15u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI254 SLI INCP net0143 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.2u l=0.06u
MI77 VDD E net110 VDD pch w=0.2u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.2u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.26u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.2u l=0.06u
MI256-M_u3 QN SLO VDD VDD pch w=0.2u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.19u l=0.06u
MI257-M_u3 net0109 SLO VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFXD1 E SE CP SI D Q QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 net0109 net108 net104 VSS nch w=0.195u l=0.06u
MI251 SLI INCPB net096 VSS nch w=0.15u l=0.06u
MI250 net096 SLO VSS VSS nch w=0.15u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI257-M_u2 net0109 SLO VSS VSS nch w=0.15u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI255-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.15u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 net0109 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI253 net0143 SLO VDD VDD pch w=0.15u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI254 SLI INCP net0143 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI257-M_u3 net0109 SLO VDD VDD pch w=0.2u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI255-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.2u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFXD2 E SE CP SI D Q QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 net0115 net108 net104 VSS nch w=0.195u l=0.06u
MI251 SLI INCPB net096 VSS nch w=0.15u l=0.06u
MI250 net096 SLO VSS VSS nch w=0.15u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI255-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI257-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI258-M_u2 net0115 SLO VSS VSS nch w=0.15u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI229-M_u2 INCPB CP VSS VSS nch w=0.195u l=0.06u
MI256-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI248-M_u2 SLO SLI VSS VSS nch w=0.195u l=0.06u
MU85-M_u2 INCP INCPB VSS VSS nch w=0.195u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 net0115 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI253 net0143 SLO VDD VDD pch w=0.15u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI254 SLI INCP net0143 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI255-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI257-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI258-M_u3 net0115 SLO VDD VDD pch w=0.2u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI229-M_u3 INCPB CP VDD VDD pch w=0.26u l=0.06u
MI256-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI248-M_u3 SLO SLI VDD VDD pch w=0.26u l=0.06u
MU85-M_u3 INCP INCPB VDD VDD pch w=0.26u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt SEDFXD4 E SE CP SI D Q QN VDD VSS
MI79 net110 E net107 VSS nch w=0.195u l=0.06u
MI135 net112 SI VSS VSS nch w=0.15u l=0.06u
MI238 net0164 INCPB VSS VSS nch w=0.2u l=0.06u
MI239 MLI d0 net0164 VSS nch w=0.2u l=0.06u
MI224 VSS E net95 VSS nch w=0.23u l=0.06u
MI222 net0116 net108 net104 VSS nch w=0.195u l=0.06u
MI251 SLI INCPB net096 VSS nch w=0.15u l=0.06u
MI250 net096 SLO VSS VSS nch w=0.15u l=0.06u
MI241 net0167 D d0 VSS nch w=0.23u l=0.06u
MI216 MLO INCP SLI VSS nch w=0.22u l=0.06u
MI119 net79 MLO VSS VSS nch w=0.15u l=0.06u
MI120 MLI INCP net79 VSS nch w=0.15u l=0.06u
MI128 net104 net147 d0 VSS nch w=0.195u l=0.06u
MI134 d0 SE net112 VSS nch w=0.15u l=0.06u
MI225 net95 net108 net0167 VSS nch w=0.23u l=0.06u
MI80 net107 net108 VSS VSS nch w=0.195u l=0.06u
MI255-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI227-M_u2 net147 E VSS VSS nch w=0.195u l=0.06u
MI257-M_u2 net0116 SLO VSS VSS nch w=0.15u l=0.06u
MI263-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI136-M_u2 net108 SE VSS VSS nch w=0.15u l=0.06u
MI264-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI265-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI259-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI266-M_u2 QN SLO VSS VSS nch w=0.39u l=0.06u
MI260-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI267-M_u2 INCPB CP VSS VSS nch w=0.31u l=0.06u
MI212-M_u2 Q SLI VSS VSS nch w=0.39u l=0.06u
MI269-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI258-M_u2 SLO SLI VSS VSS nch w=0.39u l=0.06u
MI268-M_u2 INCP INCPB VSS VSS nch w=0.25u l=0.06u
MI123-M_u2 MLO MLI VSS VSS nch w=0.35u l=0.06u
MI221 net0116 E net162 VDD pch w=0.26u l=0.06u
MI129 net162 SE d0 VDD pch w=0.26u l=0.06u
MI236 VDD INCP net0133 VDD pch w=0.27u l=0.06u
MI242 net0168 D d0 VDD pch w=0.38u l=0.06u
MI253 net0143 SLO VDD VDD pch w=0.15u l=0.06u
MI133 net177 net108 d0 VDD pch w=0.165u l=0.06u
MI226 VDD net110 net0168 VDD pch w=0.38u l=0.06u
MI254 SLI INCP net0143 VDD pch w=0.15u l=0.06u
MI210 MLO INCPB SLI VDD pch w=0.335u l=0.06u
MI235 net0133 d0 MLI VDD pch w=0.27u l=0.06u
MI102 net144 MLO VDD VDD pch w=0.15u l=0.06u
MI103 MLI INCPB net144 VDD pch w=0.15u l=0.06u
MI74 VDD net108 net110 VDD pch w=0.26u l=0.06u
MI77 VDD E net110 VDD pch w=0.26u l=0.06u
MI131 VDD SI net177 VDD pch w=0.165u l=0.06u
MI255-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI227-M_u3 net147 E VDD VDD pch w=0.25u l=0.06u
MI257-M_u3 net0116 SLO VDD VDD pch w=0.2u l=0.06u
MI263-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI136-M_u3 net108 SE VDD VDD pch w=0.2u l=0.06u
MI264-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI265-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI259-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI266-M_u3 QN SLO VDD VDD pch w=0.52u l=0.06u
MI260-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI267-M_u3 INCPB CP VDD VDD pch w=0.52u l=0.06u
MI212-M_u3 Q SLI VDD VDD pch w=0.52u l=0.06u
MI269-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
MI258-M_u3 SLO SLI VDD VDD pch w=0.5u l=0.06u
MI268-M_u3 INCP INCPB VDD VDD pch w=0.52u l=0.06u
MI123-M_u3 MLO MLI VDD VDD pch w=0.38u l=0.06u
.ends
.subckt TIEH Z VDD VSS
M_u2 net6 net6 VSS VSS nch w=0.41u l=0.06u
M_u1 Z net6 VDD VDD pch w=0.54u l=0.06u
.ends
.subckt TIEL ZN VDD VSS
M_u2 ZN net6 VSS VSS nch w=0.41u l=0.06u
M_u1 net6 net6 VDD VDD pch w=0.54u l=0.06u
.ends
.subckt XNR2D0 A1 A2 ZN VDD VSS
MI0-M_u3 net4 A1 net14 VSS nch w=0.195u l=0.06u
M_u7-M_u3 net6 net10 net14 VSS nch w=0.19u l=0.06u
M_u2-M_u2 net4 A2 VSS VSS nch w=0.195u l=0.06u
M_u5-M_u2 net6 net4 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 ZN net14 VSS VSS nch w=0.195u l=0.06u
M_u8-M_u2 net10 A1 VSS VSS nch w=0.2u l=0.06u
MI0-M_u2 net4 net10 net14 VDD pch w=0.26u l=0.06u
M_u7-M_u2 net6 A1 net14 VDD pch w=0.26u l=0.06u
M_u2-M_u3 net4 A2 VDD VDD pch w=0.26u l=0.06u
M_u5-M_u3 net6 net4 VDD VDD pch w=0.21u l=0.06u
M_u4-M_u3 ZN net14 VDD VDD pch w=0.26u l=0.06u
M_u8-M_u3 net10 A1 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR2D1 A1 A2 ZN VDD VSS
M_u2-M_u2 net4 A2 VSS VSS nch w=0.39u l=0.06u
M_u5-M_u2 net6 net4 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 ZN net14 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net10 A1 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u3 net4 A1 net14 VSS nch w=0.225u l=0.06u
MI0-M_u3 net6 net10 net14 VSS nch w=0.19u l=0.06u
M_u2-M_u3 net4 A2 VDD VDD pch w=0.52u l=0.06u
M_u5-M_u3 net6 net4 VDD VDD pch w=0.26u l=0.06u
M_u4-M_u3 ZN net14 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net10 A1 VDD VDD pch w=0.26u l=0.06u
M_u6-M_u2 net4 net10 net14 VDD pch w=0.37u l=0.06u
MI0-M_u2 net6 A1 net14 VDD pch w=0.235u l=0.06u
.ends
.subckt XNR2D2 A1 A2 ZN VDD VSS
MI1-M_u2 ZN net14 VSS VSS nch w=0.39u l=0.06u
M_u2-M_u2 net4 A2 VSS VSS nch w=0.39u l=0.06u
M_u5-M_u2 net6 net4 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 ZN net14 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net10 A1 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u3 net4 A1 net14 VSS nch w=0.225u l=0.06u
MI0-M_u3 net6 net10 net14 VSS nch w=0.19u l=0.06u
MI1-M_u3 ZN net14 VDD VDD pch w=0.52u l=0.06u
M_u2-M_u3 net4 A2 VDD VDD pch w=0.52u l=0.06u
M_u5-M_u3 net6 net4 VDD VDD pch w=0.26u l=0.06u
M_u4-M_u3 ZN net14 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net10 A1 VDD VDD pch w=0.26u l=0.06u
M_u6-M_u2 net4 net10 net14 VDD pch w=0.37u l=0.06u
MI0-M_u2 net6 A1 net14 VDD pch w=0.235u l=0.06u
.ends
.subckt XNR2D4 A1 A2 ZN VDD VSS
MI6_0-M_u3 net27 A1 net35 VSS nch w=0.3u l=0.06u
MI6_1-M_u3 net27 A1 net35 VSS nch w=0.3u l=0.06u
MI0_0-M_u3 net26 net24 net35 VSS nch w=0.31u l=0.06u
MI0_1-M_u3 net26 net24 net35 VSS nch w=0.31u l=0.06u
MI12-M_u2 net26 net27 VSS VSS nch w=0.39u l=0.06u
MI9-M_u2 ZN net35 VSS VSS nch w=0.39u l=0.06u
MI8-M_u2 ZN net35 VSS VSS nch w=0.39u l=0.06u
MI7-M_u2 ZN net35 VSS VSS nch w=0.39u l=0.06u
MI3_0-M_u2 net27 A2 VSS VSS nch w=0.39u l=0.06u
MI3_1-M_u2 net27 A2 VSS VSS nch w=0.39u l=0.06u
MI3_2-M_u2 net27 A2 VSS VSS nch w=0.39u l=0.06u
MI5-M_u2 ZN net35 VSS VSS nch w=0.39u l=0.06u
MI13-M_u2 net24 A1 VSS VSS nch w=0.29u l=0.06u
MI6_0-M_u2 net27 net24 net35 VDD pch w=0.45u l=0.06u
MI6_1-M_u2 net27 net24 net35 VDD pch w=0.45u l=0.06u
MI0_0-M_u2 net26 A1 net35 VDD pch w=0.45u l=0.06u
MI0_1-M_u2 net26 A1 net35 VDD pch w=0.45u l=0.06u
MI12-M_u3 net26 net27 VDD VDD pch w=0.52u l=0.06u
MI9-M_u3 ZN net35 VDD VDD pch w=0.52u l=0.06u
MI8-M_u3 ZN net35 VDD VDD pch w=0.52u l=0.06u
MI7-M_u3 ZN net35 VDD VDD pch w=0.52u l=0.06u
MI3_0-M_u3 net27 A2 VDD VDD pch w=0.52u l=0.06u
MI3_1-M_u3 net27 A2 VDD VDD pch w=0.52u l=0.06u
MI3_2-M_u3 net27 A2 VDD VDD pch w=0.52u l=0.06u
MI5-M_u3 ZN net35 VDD VDD pch w=0.52u l=0.06u
MI13-M_u3 net24 A1 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt XNR3D0 A1 A2 A3 ZN VDD VSS
MI8-M_u3 net11 A2 net17 VSS nch w=0.195u l=0.06u
MU11-M_u3 net5 net17 net21 VSS nch w=0.195u l=0.06u
MI5-M_u2 net5 A3 VSS VSS nch w=0.195u l=0.06u
MU22-M_u2 ZN net21 VSS VSS nch w=0.195u l=0.06u
M_u8-M_u2 net16 A2 VSS VSS nch w=0.195u l=0.06u
MI4-M_u2 net11 A1 VSS VSS nch w=0.195u l=0.06u
MI7-M_u2 net13 net17 VSS VSS nch w=0.195u l=0.06u
MI2-MU3 net17 net16 XI2-net16 VSS nch w=0.195u l=0.06u
MI2-MU4 XI2-net16 net11 VSS VSS nch w=0.195u l=0.06u
MU21-MU3 net21 net13 XU21-net16 VSS nch w=0.195u l=0.06u
MU21-MU4 XU21-net16 net5 VSS VSS nch w=0.195u l=0.06u
MI8-M_u2 net11 net16 net17 VDD pch w=0.26u l=0.06u
MU11-M_u2 net5 net13 net21 VDD pch w=0.26u l=0.06u
MI5-M_u3 net5 A3 VDD VDD pch w=0.26u l=0.06u
MU22-M_u3 ZN net21 VDD VDD pch w=0.26u l=0.06u
M_u8-M_u3 net16 A2 VDD VDD pch w=0.26u l=0.06u
MI4-M_u3 net11 A1 VDD VDD pch w=0.26u l=0.06u
MI7-M_u3 net13 net17 VDD VDD pch w=0.26u l=0.06u
MI2-MU2 net17 A2 XI2-net6 VDD pch w=0.26u l=0.06u
MI2-MU1 XI2-net6 net11 VDD VDD pch w=0.26u l=0.06u
MU21-MU2 net21 net17 XU21-net6 VDD pch w=0.26u l=0.06u
MU21-MU1 XU21-net6 net5 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR3D1 A1 A2 A3 ZN VDD VSS
M_u6-M_u3 net11 A2 net17 VSS nch w=0.195u l=0.06u
MU11-M_u3 net5 net17 net21 VSS nch w=0.28u l=0.06u
MI1-M_u2 net5 A3 VSS VSS nch w=0.39u l=0.06u
MU22-M_u2 ZN net21 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net16 A2 VSS VSS nch w=0.195u l=0.06u
M_u2-M_u2 net11 A1 VSS VSS nch w=0.39u l=0.06u
MU12-M_u2 net13 net17 VSS VSS nch w=0.195u l=0.06u
MI0-MU3 net17 net16 XI0-net16 VSS nch w=0.21u l=0.06u
MI0-MU4 XI0-net16 net11 VSS VSS nch w=0.21u l=0.06u
MI3-MU3 net21 net13 XI3-net16 VSS nch w=0.23u l=0.06u
MI3-MU4 XI3-net16 net5 VSS VSS nch w=0.23u l=0.06u
M_u6-M_u2 net11 net16 net17 VDD pch w=0.26u l=0.06u
MU11-M_u2 net5 net13 net21 VDD pch w=0.45u l=0.06u
MI1-M_u3 net5 A3 VDD VDD pch w=0.52u l=0.06u
MU22-M_u3 ZN net21 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net16 A2 VDD VDD pch w=0.26u l=0.06u
M_u2-M_u3 net11 A1 VDD VDD pch w=0.52u l=0.06u
MU12-M_u3 net13 net17 VDD VDD pch w=0.26u l=0.06u
MI0-MU2 net17 A2 XI0-net6 VDD pch w=0.36u l=0.06u
MI0-MU1 XI0-net6 net11 VDD VDD pch w=0.34u l=0.06u
MI3-MU2 net21 net17 XI3-net6 VDD pch w=0.32u l=0.06u
MI3-MU1 XI3-net6 net5 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR3D2 A1 A2 A3 ZN VDD VSS
MI8-M_u2 net42 net11 VSS VSS nch w=0.19u l=0.06u
MI5-M_u2 net44 net5 VSS VSS nch w=0.195u l=0.06u
MI7-M_u2 net5 A3 VSS VSS nch w=0.39u l=0.06u
MU22_0-M_u2 ZN net36 VSS VSS nch w=0.39u l=0.06u
MU22_1-M_u2 ZN net36 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net16 A2 VSS VSS nch w=0.195u l=0.06u
M_u2-M_u2 net11 A1 VSS VSS nch w=0.39u l=0.06u
MU12-M_u2 net54 net32 VSS VSS nch w=0.195u l=0.06u
MI3-M_u3 net42 net16 net32 VSS nch w=0.19u l=0.06u
M_u6-M_u3 net11 A2 net32 VSS nch w=0.195u l=0.06u
MU11-M_u3 net5 net32 net36 VSS nch w=0.3u l=0.06u
MI4-M_u3 net44 net54 net36 VSS nch w=0.32u l=0.06u
MI8-M_u3 net42 net11 VDD VDD pch w=0.26u l=0.06u
MI5-M_u3 net44 net5 VDD VDD pch w=0.26u l=0.06u
MI7-M_u3 net5 A3 VDD VDD pch w=0.52u l=0.06u
MU22_0-M_u3 ZN net36 VDD VDD pch w=0.52u l=0.06u
MU22_1-M_u3 ZN net36 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net16 A2 VDD VDD pch w=0.26u l=0.06u
M_u2-M_u3 net11 A1 VDD VDD pch w=0.52u l=0.06u
MU12-M_u3 net54 net32 VDD VDD pch w=0.26u l=0.06u
MI3-M_u2 net42 A2 net32 VDD pch w=0.235u l=0.06u
M_u6-M_u2 net11 net16 net32 VDD pch w=0.26u l=0.06u
MU11-M_u2 net5 net54 net36 VDD pch w=0.45u l=0.06u
MI4-M_u2 net44 net32 net36 VDD pch w=0.45u l=0.06u
.ends
.subckt XNR3D4 A1 A2 A3 ZN VDD VSS
M_u6-M_u3 net27 A2 net26 VSS nch w=0.195u l=0.06u
MI2-M_u3 net39 net25 net26 VSS nch w=0.19u l=0.06u
MU11-M_u3 p1 net26 p0 VSS nch w=0.25u l=0.06u
MI5-M_u3 net045 net40 p0 VSS nch w=0.32u l=0.06u
MI7-M_u2 net39 net27 VSS VSS nch w=0.19u l=0.06u
MI8-M_u2 net045 p1 VSS VSS nch w=0.65u l=0.06u
MI1_0-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MI1_1-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MI1_2-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MU22_0-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU22_1-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU22_2-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU22_3-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net25 A2 VSS VSS nch w=0.195u l=0.06u
M_u2_0-M_u2 net27 A1 VSS VSS nch w=0.39u l=0.06u
M_u2_1-M_u2 net27 A1 VSS VSS nch w=0.39u l=0.06u
M_u2_2-M_u2 net27 A1 VSS VSS nch w=0.39u l=0.06u
MU12-M_u2 net40 net26 VSS VSS nch w=0.39u l=0.06u
M_u6-M_u2 net27 net25 net26 VDD pch w=0.265u l=0.06u
MI2-M_u2 net39 A2 net26 VDD pch w=0.265u l=0.06u
MU11-M_u2 p1 net40 p0 VDD pch w=0.45u l=0.06u
MI5-M_u2 net045 net26 p0 VDD pch w=0.43u l=0.06u
MI7-M_u3 net39 net27 VDD VDD pch w=0.34u l=0.06u
MI8-M_u3 net045 p1 VDD VDD pch w=0.835u l=0.06u
MI1_0-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MI1_1-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MI1_2-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MU22_0-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU22_1-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU22_2-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU22_3-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net25 A2 VDD VDD pch w=0.26u l=0.06u
M_u2_0-M_u3 net27 A1 VDD VDD pch w=0.52u l=0.06u
M_u2_1-M_u3 net27 A1 VDD VDD pch w=0.52u l=0.06u
M_u2_2-M_u3 net27 A1 VDD VDD pch w=0.52u l=0.06u
MU12-M_u3 net40 net26 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt XNR4D0 A1 A2 A3 A4 ZN VDD VSS
MI21 net24 A1 net046 VSS nch w=0.195u l=0.06u
MI22 net046 net32 VSS VSS nch w=0.195u l=0.06u
MI15-M_u3 net28 net20 net64 VSS nch w=0.195u l=0.06u
MI8-M_u3 net24 net30 net32 VSS nch w=0.195u l=0.06u
MI17-M_u3 net28 net40 net24 VSS nch w=0.195u l=0.06u
MI11-M_u3 net20 A4 net108 VSS nch w=0.195u l=0.06u
MI9-M_u3 net20 net106 net104 VSS nch w=0.195u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI18-M_u2 net32 A2 VSS VSS nch w=0.195u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20-M_u2 ZN net28 VSS VSS nch w=0.195u l=0.06u
MI19-M_u2 net104 A3 VSS VSS nch w=0.195u l=0.06u
MI16-M_u2 net64 net24 VSS VSS nch w=0.195u l=0.06u
MU14-M_u2 net40 net20 VSS VSS nch w=0.195u l=0.06u
MI20 net24 net30 net045 VDD pch w=0.26u l=0.06u
M_u2 net045 net32 VDD VDD pch w=0.26u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI8-M_u2 net24 A1 net32 VDD pch w=0.26u l=0.06u
MI17-M_u2 net28 net20 net24 VDD pch w=0.26u l=0.06u
MI11-M_u2 net20 net106 net108 VDD pch w=0.26u l=0.06u
MI9-M_u2 net20 A4 net104 VDD pch w=0.26u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI18-M_u3 net32 A2 VDD VDD pch w=0.26u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20-M_u3 ZN net28 VDD VDD pch w=0.26u l=0.06u
MI19-M_u3 net104 A3 VDD VDD pch w=0.26u l=0.06u
MI16-M_u3 net64 net24 VDD VDD pch w=0.26u l=0.06u
MU14-M_u3 net40 net20 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR4D1 A1 A2 A3 A4 ZN VDD VSS
MI21 net24 A1 net043 VSS nch w=0.195u l=0.06u
MI22 net043 net32 VSS VSS nch w=0.195u l=0.06u
MI15-M_u3 net28 net20 net64 VSS nch w=0.195u l=0.06u
MI8-M_u3 net24 net30 net32 VSS nch w=0.195u l=0.06u
MI17-M_u3 net28 net40 net24 VSS nch w=0.195u l=0.06u
MI11-M_u3 net20 A4 net108 VSS nch w=0.195u l=0.06u
MI9-M_u3 net20 net106 net104 VSS nch w=0.195u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net104 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20-M_u2 ZN net28 VSS VSS nch w=0.39u l=0.06u
MI1-M_u2 net32 A2 VSS VSS nch w=0.39u l=0.06u
MI16-M_u2 net64 net24 VSS VSS nch w=0.195u l=0.06u
MU14-M_u2 net40 net20 VSS VSS nch w=0.195u l=0.06u
M_u2 net049 net32 VDD VDD pch w=0.26u l=0.06u
MI20 net24 net30 net049 VDD pch w=0.26u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI8-M_u2 net24 A1 net32 VDD pch w=0.26u l=0.06u
MI17-M_u2 net28 net20 net24 VDD pch w=0.26u l=0.06u
MI11-M_u2 net20 net106 net108 VDD pch w=0.26u l=0.06u
MI9-M_u2 net20 A4 net104 VDD pch w=0.26u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net104 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20-M_u3 ZN net28 VDD VDD pch w=0.52u l=0.06u
MI1-M_u3 net32 A2 VDD VDD pch w=0.52u l=0.06u
MI16-M_u3 net64 net24 VDD VDD pch w=0.26u l=0.06u
MU14-M_u3 net40 net20 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR4D2 A1 A2 A3 A4 ZN VDD VSS
MI15-M_u3 net28 net20 net64 VSS nch w=0.195u l=0.06u
MI8-M_u3 net24 net30 net32 VSS nch w=0.195u l=0.06u
MI6-M_u3 net24 A1 net56 VSS nch w=0.195u l=0.06u
MI17-M_u3 net28 net40 net24 VSS nch w=0.195u l=0.06u
MI11-M_u3 net20 A4 net108 VSS nch w=0.195u l=0.06u
MI9-M_u3 net20 net106 net104 VSS nch w=0.195u l=0.06u
MI19-M_u2 net56 net32 VSS VSS nch w=0.195u l=0.06u
MI21-M_u2 net64 net24 VSS VSS nch w=0.21u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net104 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20_0-M_u2 ZN net28 VSS VSS nch w=0.39u l=0.06u
MU20_1-M_u2 ZN net28 VSS VSS nch w=0.39u l=0.06u
MI1-M_u2 net32 A2 VSS VSS nch w=0.39u l=0.06u
MU14-M_u2 net40 net20 VSS VSS nch w=0.195u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI8-M_u2 net24 A1 net32 VDD pch w=0.26u l=0.06u
MI6-M_u2 net24 net30 net56 VDD pch w=0.26u l=0.06u
MI17-M_u2 net28 net20 net24 VDD pch w=0.26u l=0.06u
MI11-M_u2 net20 net106 net108 VDD pch w=0.26u l=0.06u
MI9-M_u2 net20 A4 net104 VDD pch w=0.26u l=0.06u
MI19-M_u3 net56 net32 VDD VDD pch w=0.26u l=0.06u
MI21-M_u3 net64 net24 VDD VDD pch w=0.34u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net104 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20_0-M_u3 ZN net28 VDD VDD pch w=0.52u l=0.06u
MU20_1-M_u3 ZN net28 VDD VDD pch w=0.52u l=0.06u
MI1-M_u3 net32 A2 VDD VDD pch w=0.52u l=0.06u
MU14-M_u3 net40 net20 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XNR4D4 A1 A2 A3 A4 ZN VDD VSS
MI15-M_u3 p0 net63 net78 VSS nch w=0.195u l=0.06u
MI8-M_u3 net79 net70 net67 VSS nch w=0.195u l=0.06u
MI6-M_u3 net79 A1 net66 VSS nch w=0.195u l=0.06u
MI17-M_u3 p0 net80 net79 VSS nch w=0.195u l=0.06u
MI11-M_u3 net63 A4 net72 VSS nch w=0.195u l=0.06u
MI9-M_u3 net63 net64 net68 VSS nch w=0.195u l=0.06u
MI13-M_u2 net64 A4 VSS VSS nch w=0.195u l=0.06u
MI7-M_u2 net66 net67 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net68 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net70 A1 VSS VSS nch w=0.195u l=0.06u
MI18-M_u2 net72 net68 VSS VSS nch w=0.19u l=0.06u
MU20_0-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU20_1-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU20_2-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MU20_3-M_u2 ZN p0 VSS VSS nch w=0.39u l=0.06u
MI1-M_u2 net67 A2 VSS VSS nch w=0.39u l=0.06u
MI16-M_u2 net78 net79 VSS VSS nch w=0.21u l=0.06u
MU14-M_u2 net80 net63 VSS VSS nch w=0.195u l=0.06u
MI15-M_u2 p0 net80 net78 VDD pch w=0.26u l=0.06u
MI8-M_u2 net79 A1 net67 VDD pch w=0.26u l=0.06u
MI6-M_u2 net79 net70 net66 VDD pch w=0.26u l=0.06u
MI17-M_u2 p0 net63 net79 VDD pch w=0.26u l=0.06u
MI11-M_u2 net63 net64 net72 VDD pch w=0.26u l=0.06u
MI9-M_u2 net63 A4 net68 VDD pch w=0.26u l=0.06u
MI13-M_u3 net64 A4 VDD VDD pch w=0.26u l=0.06u
MI7-M_u3 net66 net67 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net68 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net70 A1 VDD VDD pch w=0.26u l=0.06u
MI18-M_u3 net72 net68 VDD VDD pch w=0.21u l=0.06u
MU20_0-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU20_1-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU20_2-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MU20_3-M_u3 ZN p0 VDD VDD pch w=0.52u l=0.06u
MI1-M_u3 net67 A2 VDD VDD pch w=0.52u l=0.06u
MI16-M_u3 net78 net79 VDD VDD pch w=0.34u l=0.06u
MU14-M_u3 net80 net63 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR2D0 A1 A2 Z VDD VSS
M_u6-M_u3 net4 net10 net14 VSS nch w=0.195u l=0.06u
MI5-M_u3 net6 A1 net14 VSS nch w=0.195u l=0.06u
MI1-M_u2 net4 A2 VSS VSS nch w=0.195u l=0.06u
M_u5-M_u2 net6 net4 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 Z net14 VSS VSS nch w=0.195u l=0.06u
MI4-M_u2 net10 A1 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u2 net4 A1 net14 VDD pch w=0.26u l=0.06u
MI5-M_u2 net6 net10 net14 VDD pch w=0.26u l=0.06u
MI1-M_u3 net4 A2 VDD VDD pch w=0.26u l=0.06u
M_u5-M_u3 net6 net4 VDD VDD pch w=0.21u l=0.06u
M_u4-M_u3 Z net14 VDD VDD pch w=0.26u l=0.06u
MI4-M_u3 net10 A1 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR2D1 A1 A2 Z VDD VSS
M_u6-M_u3 net4 net10 net14 VSS nch w=0.32u l=0.06u
MI1-M_u3 net6 A1 net14 VSS nch w=0.31u l=0.06u
M_u2-M_u2 net4 A2 VSS VSS nch w=0.39u l=0.06u
M_u5-M_u2 net6 net4 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 Z net14 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net10 A1 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u2 net4 A1 net14 VDD pch w=0.34u l=0.06u
MI1-M_u2 net6 net10 net14 VDD pch w=0.31u l=0.06u
M_u2-M_u3 net4 A2 VDD VDD pch w=0.52u l=0.06u
M_u5-M_u3 net6 net4 VDD VDD pch w=0.21u l=0.06u
M_u4-M_u3 Z net14 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net10 A1 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR2D2 A1 A2 Z VDD VSS
MI2-M_u2 Z net27 VSS VSS nch w=0.39u l=0.06u
M_u2-M_u2 net23 A2 VSS VSS nch w=0.39u l=0.06u
M_u5-M_u2 net21 net23 VSS VSS nch w=0.19u l=0.06u
M_u4-M_u2 Z net27 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net17 A1 VSS VSS nch w=0.195u l=0.06u
MI1-M_u3 net21 A1 net27 VSS nch w=0.31u l=0.06u
M_u6-M_u3 net23 net17 net27 VSS nch w=0.32u l=0.06u
MI2-M_u3 Z net27 VDD VDD pch w=0.52u l=0.06u
M_u2-M_u3 net23 A2 VDD VDD pch w=0.52u l=0.06u
M_u5-M_u3 net21 net23 VDD VDD pch w=0.26u l=0.06u
M_u4-M_u3 Z net27 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net17 A1 VDD VDD pch w=0.26u l=0.06u
MI1-M_u2 net21 net17 net27 VDD pch w=0.31u l=0.06u
M_u6-M_u2 net23 A1 net27 VDD pch w=0.34u l=0.06u
.ends
.subckt XOR2D4 A1 A2 Z VDD VSS
MI3_0-M_u3 net026 net29 p0 VSS nch w=0.3u l=0.06u
MI3_1-M_u3 net026 net29 p0 VSS nch w=0.3u l=0.06u
MI4_0-M_u3 net6 A1 p0 VSS nch w=0.31u l=0.06u
MI4_1-M_u3 net6 A1 p0 VSS nch w=0.31u l=0.06u
M_u2_0-M_u2 net026 A2 VSS VSS nch w=0.39u l=0.06u
M_u2_1-M_u2 net026 A2 VSS VSS nch w=0.39u l=0.06u
M_u2_2-M_u2 net026 A2 VSS VSS nch w=0.39u l=0.06u
M_u5-M_u2 net6 net026 VSS VSS nch w=0.39u l=0.06u
M_u4_0-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_1-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_2-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u4_3-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net29 A1 VSS VSS nch w=0.39u l=0.06u
MI3_0-M_u2 net026 A1 p0 VDD pch w=0.45u l=0.06u
MI3_1-M_u2 net026 A1 p0 VDD pch w=0.45u l=0.06u
MI4_0-M_u2 net6 net29 p0 VDD pch w=0.45u l=0.06u
MI4_1-M_u2 net6 net29 p0 VDD pch w=0.45u l=0.06u
M_u2_0-M_u3 net026 A2 VDD VDD pch w=0.52u l=0.06u
M_u2_1-M_u3 net026 A2 VDD VDD pch w=0.52u l=0.06u
M_u2_2-M_u3 net026 A2 VDD VDD pch w=0.52u l=0.06u
M_u5-M_u3 net6 net026 VDD VDD pch w=0.52u l=0.06u
M_u4_0-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u4_1-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u4_2-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u4_3-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net29 A1 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt XOR3D0 A1 A2 A3 Z VDD VSS
M_u6-M_u3 net19 net17 net25 VSS nch w=0.195u l=0.06u
MU18-M_u3 net13 net25 net29 VSS nch w=0.195u l=0.06u
MI1-M_u2 Z net29 VSS VSS nch w=0.195u l=0.06u
MI3-M_u2 net13 A3 VSS VSS nch w=0.195u l=0.06u
MI7-M_u2 net17 A2 VSS VSS nch w=0.195u l=0.06u
MI2-M_u2 net19 A1 VSS VSS nch w=0.195u l=0.06u
MI6-M_u2 net21 net25 VSS VSS nch w=0.195u l=0.06u
MU33-MU3 net29 net21 XU33-net16 VSS nch w=0.195u l=0.06u
MU33-MU4 XU33-net16 net13 VSS VSS nch w=0.195u l=0.06u
MI5-MU3 net25 A2 XI5-net16 VSS nch w=0.195u l=0.06u
MI5-MU4 XI5-net16 net19 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u2 net19 A2 net25 VDD pch w=0.26u l=0.06u
MU18-M_u2 net13 net21 net29 VDD pch w=0.26u l=0.06u
MI1-M_u3 Z net29 VDD VDD pch w=0.26u l=0.06u
MI3-M_u3 net13 A3 VDD VDD pch w=0.26u l=0.06u
MI7-M_u3 net17 A2 VDD VDD pch w=0.26u l=0.06u
MI2-M_u3 net19 A1 VDD VDD pch w=0.26u l=0.06u
MI6-M_u3 net21 net25 VDD VDD pch w=0.26u l=0.06u
MU33-MU2 net29 net25 XU33-net6 VDD pch w=0.26u l=0.06u
MU33-MU1 XU33-net6 net13 VDD VDD pch w=0.26u l=0.06u
MI5-MU2 net25 net17 XI5-net6 VDD pch w=0.26u l=0.06u
MI5-MU1 XI5-net6 net19 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR3D1 A1 A2 A3 Z VDD VSS
M_u6-M_u3 net19 net17 net25 VSS nch w=0.195u l=0.06u
MU18-M_u3 net13 net25 net29 VSS nch w=0.28u l=0.06u
MU13-M_u2 net13 A3 VSS VSS nch w=0.39u l=0.06u
MU14-M_u2 Z net29 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net17 A2 VSS VSS nch w=0.195u l=0.06u
M_u2-M_u2 net19 A1 VSS VSS nch w=0.39u l=0.06u
M_u4-M_u2 net21 net25 VSS VSS nch w=0.195u l=0.06u
MU33-MU3 net29 net21 XU33-net16 VSS nch w=0.23u l=0.06u
MU33-MU4 XU33-net16 net13 VSS VSS nch w=0.23u l=0.06u
MI0-MU3 net25 A2 XI0-net16 VSS nch w=0.195u l=0.06u
MI0-MU4 XI0-net16 net19 VSS VSS nch w=0.195u l=0.06u
M_u6-M_u2 net19 A2 net25 VDD pch w=0.26u l=0.06u
MU18-M_u2 net13 net21 net29 VDD pch w=0.45u l=0.06u
MU13-M_u3 net13 A3 VDD VDD pch w=0.52u l=0.06u
MU14-M_u3 Z net29 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net17 A2 VDD VDD pch w=0.26u l=0.06u
M_u2-M_u3 net19 A1 VDD VDD pch w=0.52u l=0.06u
M_u4-M_u3 net21 net25 VDD VDD pch w=0.26u l=0.06u
MU33-MU2 net29 net25 XU33-net6 VDD pch w=0.32u l=0.06u
MU33-MU1 XU33-net6 net13 VDD VDD pch w=0.26u l=0.06u
MI0-MU2 net25 net17 XI0-net6 VDD pch w=0.26u l=0.06u
MI0-MU1 XI0-net6 net19 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR3D2 A1 A2 A3 Z VDD VSS
MI6-M_u2 net13 A3 VSS VSS nch w=0.39u l=0.06u
MI8-M_u2 net44 net19 VSS VSS nch w=0.19u l=0.06u
MI9-M_u2 net42 net13 VSS VSS nch w=0.15u l=0.06u
MU14_0-M_u2 Z net32 VSS VSS nch w=0.39u l=0.06u
MU14_1-M_u2 Z net32 VSS VSS nch w=0.39u l=0.06u
MI7-M_u2 net17 A2 VSS VSS nch w=0.195u l=0.06u
M_u2-M_u2 net19 A1 VSS VSS nch w=0.39u l=0.06u
M_u4-M_u2 net21 net25 VSS VSS nch w=0.195u l=0.06u
MI3-M_u3 net42 net21 net32 VSS nch w=0.19u l=0.06u
M_u6-M_u3 net19 net17 net25 VSS nch w=0.195u l=0.06u
MI1-M_u3 net44 A2 net25 VSS nch w=0.195u l=0.06u
MU18-M_u3 net13 net25 net32 VSS nch w=0.27u l=0.06u
MI6-M_u3 net13 A3 VDD VDD pch w=0.52u l=0.06u
MI8-M_u3 net44 net19 VDD VDD pch w=0.21u l=0.06u
MI9-M_u3 net42 net13 VDD VDD pch w=0.24u l=0.06u
MU14_0-M_u3 Z net32 VDD VDD pch w=0.52u l=0.06u
MU14_1-M_u3 Z net32 VDD VDD pch w=0.52u l=0.06u
MI7-M_u3 net17 A2 VDD VDD pch w=0.26u l=0.06u
M_u2-M_u3 net19 A1 VDD VDD pch w=0.52u l=0.06u
M_u4-M_u3 net21 net25 VDD VDD pch w=0.24u l=0.06u
MI3-M_u2 net42 net25 net32 VDD pch w=0.33u l=0.06u
M_u6-M_u2 net19 A2 net25 VDD pch w=0.26u l=0.06u
MI1-M_u2 net44 net17 net25 VDD pch w=0.26u l=0.06u
MU18-M_u2 net13 net21 net32 VDD pch w=0.45u l=0.06u
.ends
.subckt XOR3D4 A1 A2 A3 Z VDD VSS
MI9-M_u3 net031 net21 p0 VSS nch w=0.32u l=0.06u
M_u6-M_u3 net29 net17 net28 VSS nch w=0.195u l=0.06u
MI1-M_u3 net28 A2 net39 VSS nch w=0.195u l=0.06u
MU18-M_u3 p1 net28 p0 VSS nch w=0.25u l=0.06u
MI7-M_u2 net39 net29 VSS VSS nch w=0.19u l=0.06u
MI8_0-M_u2 net031 p1 VSS VSS nch w=0.39u l=0.06u
MI8_1-M_u2 net031 p1 VSS VSS nch w=0.39u l=0.06u
MU13_0-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MU13_1-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MU13_2-M_u2 p1 A3 VSS VSS nch w=0.39u l=0.06u
MU14_0-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU14_1-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU14_2-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU14_3-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI11-M_u2 net17 A2 VSS VSS nch w=0.195u l=0.06u
M_u2_0-M_u2 net29 A1 VSS VSS nch w=0.39u l=0.06u
M_u2_1-M_u2 net29 A1 VSS VSS nch w=0.39u l=0.06u
M_u2_2-M_u2 net29 A1 VSS VSS nch w=0.39u l=0.06u
M_u4-M_u2 net21 net28 VSS VSS nch w=0.39u l=0.06u
MI9-M_u2 net031 net28 p0 VDD pch w=0.45u l=0.06u
M_u6-M_u2 net29 A2 net28 VDD pch w=0.26u l=0.06u
MI1-M_u2 net28 net17 net39 VDD pch w=0.26u l=0.06u
MU18-M_u2 p1 net21 p0 VDD pch w=0.45u l=0.06u
MI7-M_u3 net39 net29 VDD VDD pch w=0.21u l=0.06u
MI8_0-M_u3 net031 p1 VDD VDD pch w=0.43u l=0.06u
MI8_1-M_u3 net031 p1 VDD VDD pch w=0.43u l=0.06u
MU13_0-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MU13_1-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MU13_2-M_u3 p1 A3 VDD VDD pch w=0.52u l=0.06u
MU14_0-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU14_1-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU14_2-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU14_3-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MI11-M_u3 net17 A2 VDD VDD pch w=0.26u l=0.06u
M_u2_0-M_u3 net29 A1 VDD VDD pch w=0.52u l=0.06u
M_u2_1-M_u3 net29 A1 VDD VDD pch w=0.52u l=0.06u
M_u2_2-M_u3 net29 A1 VDD VDD pch w=0.52u l=0.06u
M_u4-M_u3 net21 net28 VDD VDD pch w=0.54u l=0.06u
.ends
.subckt XOR4D0 A1 A2 A3 A4 Z VDD VSS
MI21 net24 A1 net050 VSS nch w=0.195u l=0.06u
MI22 net050 net32 VSS VSS nch w=0.195u l=0.06u
MI15-M_u3 net28 net20 net64 VSS nch w=0.195u l=0.06u
MI8-M_u3 net24 net30 net32 VSS nch w=0.195u l=0.06u
MI17-M_u3 net28 net40 net24 VSS nch w=0.195u l=0.06u
MI11-M_u3 net40 A4 net108 VSS nch w=0.195u l=0.06u
MI9-M_u3 net40 net106 net104 VSS nch w=0.195u l=0.06u
MI19-M_u2 net20 net40 VSS VSS nch w=0.195u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net104 A3 VSS VSS nch w=0.195u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20-M_u2 Z net28 VSS VSS nch w=0.195u l=0.06u
MI1-M_u2 net32 A2 VSS VSS nch w=0.195u l=0.06u
MI16-M_u2 net64 net24 VSS VSS nch w=0.195u l=0.06u
MI20 net24 net30 net045 VDD pch w=0.26u l=0.06u
M_u2 net045 net32 VDD VDD pch w=0.26u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI8-M_u2 net24 A1 net32 VDD pch w=0.26u l=0.06u
MI17-M_u2 net28 net20 net24 VDD pch w=0.26u l=0.06u
MI11-M_u2 net40 net106 net108 VDD pch w=0.26u l=0.06u
MI9-M_u2 net40 A4 net104 VDD pch w=0.26u l=0.06u
MI19-M_u3 net20 net40 VDD VDD pch w=0.26u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net104 A3 VDD VDD pch w=0.26u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20-M_u3 Z net28 VDD VDD pch w=0.26u l=0.06u
MI1-M_u3 net32 A2 VDD VDD pch w=0.26u l=0.06u
MI16-M_u3 net64 net24 VDD VDD pch w=0.26u l=0.06u
.ends
.subckt XOR4D1 A1 A2 A3 A4 Z VDD VSS
MI21 net24 A1 net048 VSS nch w=0.195u l=0.06u
MI29 net048 net32 VSS VSS nch w=0.195u l=0.06u
MI15-M_u3 net28 net20 net64 VSS nch w=0.21u l=0.06u
MI26-M_u3 net24 net30 net32 VSS nch w=0.32u l=0.06u
MI28-M_u3 net40 net106 net104 VSS nch w=0.32u l=0.06u
MI27-M_u3 net40 A4 net108 VSS nch w=0.29u l=0.06u
MI24-M_u3 net28 net40 net24 VSS nch w=0.295u l=0.06u
MI22-M_u2 net64 net24 VSS VSS nch w=0.21u l=0.06u
MI23-M_u2 net20 net40 VSS VSS nch w=0.39u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net104 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20-M_u2 Z net28 VSS VSS nch w=0.39u l=0.06u
MI1-M_u2 net32 A2 VSS VSS nch w=0.39u l=0.06u
MI20 net24 net30 net043 VDD pch w=0.26u l=0.06u
M_u2 net043 net32 VDD VDD pch w=0.26u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI26-M_u2 net24 A1 net32 VDD pch w=0.415u l=0.06u
MI28-M_u2 net40 A4 net104 VDD pch w=0.32u l=0.06u
MI27-M_u2 net40 net106 net108 VDD pch w=0.32u l=0.06u
MI24-M_u2 net28 net20 net24 VDD pch w=0.45u l=0.06u
MI22-M_u3 net64 net24 VDD VDD pch w=0.34u l=0.06u
MI23-M_u3 net20 net40 VDD VDD pch w=0.37u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net104 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20-M_u3 Z net28 VDD VDD pch w=0.52u l=0.06u
MI1-M_u3 net32 A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt XOR4D2 A1 A2 A3 A4 Z VDD VSS
MI15-M_u3 net28 net20 net64 VSS nch w=0.21u l=0.06u
MI26-M_u3 net24 net30 net32 VSS nch w=0.32u l=0.06u
MI28-M_u3 net40 net106 net104 VSS nch w=0.32u l=0.06u
MI27-M_u3 net40 A4 net108 VSS nch w=0.29u l=0.06u
MI24-M_u3 net28 net40 net24 VSS nch w=0.295u l=0.06u
MI25-M_u3 net24 A1 net56 VSS nch w=0.195u l=0.06u
MI22-M_u2 net64 net24 VSS VSS nch w=0.21u l=0.06u
MI29-M_u2 Z net28 VSS VSS nch w=0.39u l=0.06u
MI23-M_u2 net20 net40 VSS VSS nch w=0.39u l=0.06u
MI13-M_u2 net106 A4 VSS VSS nch w=0.195u l=0.06u
MI7-M_u2 net56 net32 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net104 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net30 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net108 net104 VSS VSS nch w=0.19u l=0.06u
MU20-M_u2 Z net28 VSS VSS nch w=0.39u l=0.06u
MI1-M_u2 net32 A2 VSS VSS nch w=0.39u l=0.06u
MI15-M_u2 net28 net40 net64 VDD pch w=0.26u l=0.06u
MI26-M_u2 net24 A1 net32 VDD pch w=0.415u l=0.06u
MI28-M_u2 net40 A4 net104 VDD pch w=0.32u l=0.06u
MI27-M_u2 net40 net106 net108 VDD pch w=0.32u l=0.06u
MI24-M_u2 net28 net20 net24 VDD pch w=0.45u l=0.06u
MI25-M_u2 net24 net30 net56 VDD pch w=0.26u l=0.06u
MI22-M_u3 net64 net24 VDD VDD pch w=0.34u l=0.06u
MI29-M_u3 Z net28 VDD VDD pch w=0.52u l=0.06u
MI23-M_u3 net20 net40 VDD VDD pch w=0.37u l=0.06u
MI13-M_u3 net106 A4 VDD VDD pch w=0.26u l=0.06u
MI7-M_u3 net56 net32 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net104 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net30 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net108 net104 VDD VDD pch w=0.21u l=0.06u
MU20-M_u3 Z net28 VDD VDD pch w=0.52u l=0.06u
MI1-M_u3 net32 A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt XOR4D4 A1 A2 A3 A4 Z VDD VSS
MI23-M_u3 net64 A1 net47 VSS nch w=0.275u l=0.06u
MI35-M_u3 net81 net66 p0 VSS nch w=0.32u l=0.06u
MI36-M_u3 net47 net63 p0 VSS nch w=0.195u l=0.06u
MI33-M_u3 net74 A4 net63 VSS nch w=0.29u l=0.06u
MI34-M_u3 net70 net68 net63 VSS nch w=0.32u l=0.06u
MI32-M_u3 net65 net72 net47 VSS nch w=0.32u l=0.06u
MI27-M_u2 net64 net65 VSS VSS nch w=0.21u l=0.06u
MI31_0-M_u2 net81 net47 VSS VSS nch w=0.39u l=0.06u
MI31_1-M_u2 net81 net47 VSS VSS nch w=0.39u l=0.06u
MI26-M_u2 net66 net63 VSS VSS nch w=0.195u l=0.06u
MI13-M_u2 net68 A4 VSS VSS nch w=0.195u l=0.06u
MI14-M_u2 net70 A3 VSS VSS nch w=0.39u l=0.06u
M_u8-M_u2 net72 A1 VSS VSS nch w=0.195u l=0.06u
MI12-M_u2 net74 net70 VSS VSS nch w=0.19u l=0.06u
MU20_0-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU20_1-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU20_2-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MU20_3-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI1_0-M_u2 net65 A2 VSS VSS nch w=0.39u l=0.06u
MI1_1-M_u2 net65 A2 VSS VSS nch w=0.39u l=0.06u
MI23-M_u2 net64 net72 net47 VDD pch w=0.26u l=0.06u
MI35-M_u2 net81 net63 p0 VDD pch w=0.42u l=0.06u
MI36-M_u2 net47 net66 p0 VDD pch w=0.24u l=0.06u
MI33-M_u2 net74 net68 net63 VDD pch w=0.32u l=0.06u
MI34-M_u2 net70 A4 net63 VDD pch w=0.32u l=0.06u
MI32-M_u2 net65 A1 net47 VDD pch w=0.335u l=0.06u
MI27-M_u3 net64 net65 VDD VDD pch w=0.34u l=0.06u
MI31_0-M_u3 net81 net47 VDD VDD pch w=0.52u l=0.06u
MI31_1-M_u3 net81 net47 VDD VDD pch w=0.52u l=0.06u
MI26-M_u3 net66 net63 VDD VDD pch w=0.26u l=0.06u
MI13-M_u3 net68 A4 VDD VDD pch w=0.26u l=0.06u
MI14-M_u3 net70 A3 VDD VDD pch w=0.52u l=0.06u
M_u8-M_u3 net72 A1 VDD VDD pch w=0.26u l=0.06u
MI12-M_u3 net74 net70 VDD VDD pch w=0.21u l=0.06u
MU20_0-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU20_1-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU20_2-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MU20_3-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
MI1_0-M_u3 net65 A2 VDD VDD pch w=0.52u l=0.06u
MI1_1-M_u3 net65 A2 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ISOHID1 ISO I Z VDD VSS
MI3-M_u2 Z net15 VSS VSS nch w=0.39u l=0.06u
MI1-M_u4 net15 I VSS VSS nch w=0.39u l=0.06u
MI1-M_u3 net15 ISO VSS VSS nch w=0.39u l=0.06u
MI3-M_u3 Z net15 VDD VDD pch w=0.52u l=0.06u
MI1-M_u1 XI1-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1-M_u2 net15 I XI1-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt ISOHID2 ISO I Z VDD VSS
MI3_0-M_u2 Z net11 VSS VSS nch w=0.39u l=0.06u
MI3_1-M_u2 Z net11 VSS VSS nch w=0.39u l=0.06u
MI1-M_u4 net11 I VSS VSS nch w=0.39u l=0.06u
MI1-M_u3 net11 ISO VSS VSS nch w=0.39u l=0.06u
MI3_0-M_u3 Z net11 VDD VDD pch w=0.52u l=0.06u
MI3_1-M_u3 Z net11 VDD VDD pch w=0.52u l=0.06u
MI1-M_u1 XI1-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1-M_u2 net11 I XI1-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt ISOHID4 ISO I Z VDD VSS
MI3_0-M_u2 Z net20 VSS VSS nch w=0.39u l=0.06u
MI3_1-M_u2 Z net20 VSS VSS nch w=0.39u l=0.06u
MI3_2-M_u2 Z net20 VSS VSS nch w=0.39u l=0.06u
MI3_3-M_u2 Z net20 VSS VSS nch w=0.39u l=0.06u
MI1-M_u4 net20 I VSS VSS nch w=0.39u l=0.06u
MI1-M_u3 net20 ISO VSS VSS nch w=0.39u l=0.06u
MI3_0-M_u3 Z net20 VDD VDD pch w=0.52u l=0.06u
MI3_1-M_u3 Z net20 VDD VDD pch w=0.52u l=0.06u
MI3_2-M_u3 Z net20 VDD VDD pch w=0.52u l=0.06u
MI3_3-M_u3 Z net20 VDD VDD pch w=0.52u l=0.06u
MI1-M_u1 XI1-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1-M_u2 net20 I XI1-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt ISOHID8 ISO I Z VDD VSS
MI3_0-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_1-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_2-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_3-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_4-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_5-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_6-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI3_7-M_u2 Z P0 VSS VSS nch w=0.39u l=0.06u
MI1_0-M_u4 P0 I VSS VSS nch w=0.39u l=0.06u
MI1_0-M_u3 P0 ISO VSS VSS nch w=0.39u l=0.06u
MI1_1-M_u4 P0 I VSS VSS nch w=0.39u l=0.06u
MI1_1-M_u3 P0 ISO VSS VSS nch w=0.39u l=0.06u
MI1_2-M_u4 P0 I VSS VSS nch w=0.39u l=0.06u
MI1_2-M_u3 P0 ISO VSS VSS nch w=0.39u l=0.06u
MI3_0-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_1-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_2-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_3-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_4-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_5-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_6-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI3_7-M_u3 Z P0 VDD VDD pch w=0.52u l=0.06u
MI1_0-M_u1 XI1_0-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1_0-M_u2 P0 I XI1_0-net8 VDD pch w=0.52u l=0.06u
MI1_1-M_u1 XI1_1-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1_1-M_u2 P0 I XI1_1-net8 VDD pch w=0.52u l=0.06u
MI1_2-M_u1 XI1_2-net8 ISO VDD VDD pch w=0.52u l=0.06u
MI1_2-M_u2 P0 I XI1_2-net8 VDD pch w=0.52u l=0.06u
.ends
.subckt ISOLOD1 ISO I Z VDD VSS
MI3-M_u3 Z net025 VDD VDD pch w=0.52u l=0.06u
MI2-M_u3 net13 ISO VDD VDD pch w=0.26u l=0.06u
M_u16 VDD net13 net025 VDD pch w=0.52u l=0.06u
MI11 VDD I net025 VDD pch w=0.52u l=0.06u
MI3-M_u2 Z net025 VSS VSS nch w=0.39u l=0.06u
MI2-M_u2 net13 ISO VSS VSS nch w=0.195u l=0.06u
MI13 net16 net13 VSS VSS nch w=0.39u l=0.06u
MI12 net025 I net16 VSS nch w=0.39u l=0.06u
.ends
.subckt ISOLOD2 ISO I Z VDD VSS
MI4 net22 net017 VSS VSS nch w=0.39u l=0.06u
MI12 net037 I net22 VSS nch w=0.39u l=0.06u
MI13-M_u2 net017 ISO VSS VSS nch w=0.195u l=0.06u
M_u3-M_u2 Z net037 VSS VSS nch w=0.39u l=0.06u
MI14-M_u2 Z net037 VSS VSS nch w=0.39u l=0.06u
M_u16 VDD net017 net037 VDD pch w=0.52u l=0.06u
MI3 VDD I net037 VDD pch w=0.52u l=0.06u
MI13-M_u3 net017 ISO VDD VDD pch w=0.26u l=0.06u
M_u3-M_u3 Z net037 VDD VDD pch w=0.52u l=0.06u
MI14-M_u3 Z net037 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt ISOLOD4 ISO I Z VDD VSS
MI13 net021 p0 VSS VSS nch w=0.39u l=0.06u
MI12 net016 I net021 VSS nch w=0.39u l=0.06u
MI4_0-M_u2 Z net016 VSS VSS nch w=0.39u l=0.06u
MI4_1-M_u2 Z net016 VSS VSS nch w=0.39u l=0.06u
MI4_2-M_u2 Z net016 VSS VSS nch w=0.39u l=0.06u
MI4_3-M_u2 Z net016 VSS VSS nch w=0.39u l=0.06u
MI2-M_u2 p0 ISO VSS VSS nch w=0.195u l=0.06u
M_u16 VDD p0 net016 VDD pch w=0.52u l=0.06u
MI11 VDD I net016 VDD pch w=0.52u l=0.06u
MI4_0-M_u3 Z net016 VDD VDD pch w=0.52u l=0.06u
MI4_1-M_u3 Z net016 VDD VDD pch w=0.52u l=0.06u
MI4_2-M_u3 Z net016 VDD VDD pch w=0.52u l=0.06u
MI4_3-M_u3 Z net016 VDD VDD pch w=0.52u l=0.06u
MI2-M_u3 p0 ISO VDD VDD pch w=0.26u l=0.06u
.ends
.subckt ISOLOD8 ISO I Z VDD VSS
MI13_0 net21<0> p0 VSS VSS nch w=0.39u l=0.06u
MI13_1 net21<1> p0 VSS VSS nch w=0.39u l=0.06u
MI13_2 net21<2> p0 VSS VSS nch w=0.39u l=0.06u
MI12_0 P1 I net21<0> VSS nch w=0.39u l=0.06u
MI12_1 P1 I net21<1> VSS nch w=0.39u l=0.06u
MI12_2 P1 I net21<2> VSS nch w=0.39u l=0.06u
MI4_0-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_1-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_2-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_3-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_4-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_5-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_6-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI4_7-M_u2 Z P1 VSS VSS nch w=0.39u l=0.06u
MI2-M_u2 p0 ISO VSS VSS nch w=0.39u l=0.06u
M_u16_0 VDD p0 P1 VDD pch w=0.52u l=0.06u
M_u16_1 VDD p0 P1 VDD pch w=0.52u l=0.06u
M_u16_2 VDD p0 P1 VDD pch w=0.52u l=0.06u
MI11_0 VDD I P1 VDD pch w=0.52u l=0.06u
MI11_1 VDD I P1 VDD pch w=0.52u l=0.06u
MI11_2 VDD I P1 VDD pch w=0.52u l=0.06u
MI4_0-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_1-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_2-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_3-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_4-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_5-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_6-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI4_7-M_u3 Z P1 VDD VDD pch w=0.52u l=0.06u
MI2-M_u3 p0 ISO VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLHLD1 I Z VDD VSS
MI1-M_u2 Z net6 VSS VSS nch w=0.39u l=0.06u
MI2-M_u2 net6 I VSS VSS nch w=0.195u l=0.06u
MI1-M_u3 Z net6 VDD VDD pch w=0.52u l=0.06u
MI2-M_u3 net6 I VDD VDD pch w=0.26u l=0.06u
.ends
.subckt LVLHLD2 I Z VDD VSS
M_u2-M_u2 net8 I VSS VSS nch w=0.39u l=0.06u
M_u3_0-M_u2 Z net8 VSS VSS nch w=0.39u l=0.06u
M_u3_1-M_u2 Z net8 VSS VSS nch w=0.39u l=0.06u
M_u2-M_u3 net8 I VDD VDD pch w=0.52u l=0.06u
M_u3_0-M_u3 Z net8 VDD VDD pch w=0.52u l=0.06u
M_u3_1-M_u3 Z net8 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLHLD4 I Z VDD VSS
M_u3_0-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u3_1-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u3_2-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u3_3-M_u2 Z p0 VSS VSS nch w=0.39u l=0.06u
M_u2_0-M_u2 p0 I VSS VSS nch w=0.39u l=0.06u
M_u2_1-M_u2 p0 I VSS VSS nch w=0.39u l=0.06u
M_u3_0-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u3_1-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u3_2-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u3_3-M_u3 Z p0 VDD VDD pch w=0.52u l=0.06u
M_u2_0-M_u3 p0 I VDD VDD pch w=0.52u l=0.06u
M_u2_1-M_u3 p0 I VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLHLD8 I Z VDD VSS
M_u2_0-M_u2 n0 I VSS VSS nch w=0.39u l=0.06u
M_u2_1-M_u2 n0 I VSS VSS nch w=0.39u l=0.06u
M_u2_2-M_u2 n0 I VSS VSS nch w=0.39u l=0.06u
M_u7_0-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_1-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_2-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_3-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_4-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_5-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_6-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u7_7-M_u2 Z n0 VSS VSS nch w=0.39u l=0.06u
M_u2_0-M_u3 n0 I VDD VDD pch w=0.52u l=0.06u
M_u2_1-M_u3 n0 I VDD VDD pch w=0.52u l=0.06u
M_u2_2-M_u3 n0 I VDD VDD pch w=0.52u l=0.06u
M_u7_0-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_1-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_2-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_3-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_4-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_5-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_6-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
M_u7_7-M_u3 Z n0 VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLLHCD1 I NSLEEP Z VDD VDDL VSS
MI16 Z net031 vvss VSS nch w=0.39u l=0.06u
MI44 net024 I vvss VSS nch w=0.39u l=0.06u
MI43_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI43_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI43_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40_0 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_1 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_2 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_3 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI42_0 net031 I vvss VSS nch w=0.39u l=0.06u
MI42_1 net031 I vvss VSS nch w=0.39u l=0.06u
MI42_2 net031 I vvss VSS nch w=0.39u l=0.06u
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net031 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net031 net34 VDD pch w=0.15u l=0.06u
MI15 VDD net031 Z VDD pch w=0.52u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.15u l=0.06u
.ends
.subckt LVLLHCD2 I NSLEEP Z VDD VDDL VSS
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net043 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net043 net34 VDD pch w=0.15u l=0.06u
MI15_0 VDD net043 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net043 Z VDD pch w=0.52u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.34u l=0.06u
MI16_0 Z net043 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net043 vvss VSS nch w=0.39u l=0.06u
MI45 net024 I vvss VSS nch w=0.39u l=0.06u
MI44_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI44_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI44_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40_0 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_1 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_2 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_3 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI43_0 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_1 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_2 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_3 net043 I vvss VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHCD4 I NSLEEP Z VDD VDDL VSS
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net038 net34 VDD VDD pch w=0.15u l=0.06u
MI15_0 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD net038 Z VDD pch w=0.52u l=0.06u
MI37 VDD net038 net34 VDD pch w=0.15u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
MI45_0 net038 I vvss VSS nch w=0.39u l=0.06u
MI45_1 net038 I vvss VSS nch w=0.39u l=0.06u
MI45_2 net038 I vvss VSS nch w=0.39u l=0.06u
MI46_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40 vvss NSLEEP VSS VSS nch w=3.11u l=0.06u
MI16_0 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_2 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_3 Z net038 vvss VSS nch w=0.39u l=0.06u
MI47 net024 I vvss VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHCD8 I NSLEEP Z VDD VDDL VSS
MI45_0 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_1 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_2 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_3 net087 I vvss VSS nch w=0.39u l=0.06u
MI46_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI16_0 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_2 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_3 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_4 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_5 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_6 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_7 Z net087 vvss VSS nch w=0.39u l=0.06u
MI40 vvss NSLEEP VSS VSS nch w=6.26u l=0.06u
MI47 net024 I vvss VSS nch w=0.39u l=0.06u
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net087 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net087 net34 VDD pch w=0.15u l=0.06u
MI15_0 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_4 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_5 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_6 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_7 VDD net087 Z VDD pch w=0.52u l=0.06u
MI41_0 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
MI41_1 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLLHD1 I Z VDD VDDL VSS
MI15 VDD net25 Z VDD pch w=0.52u l=0.06u
MI5 VDD net25 net34 VDD pch w=0.15u l=0.06u
MI19 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI17 net25 net34 VDD VDD pch w=0.15u l=0.06u
MI6_0 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_1 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_2 net25 I VSS VSS nch w=0.39u l=0.06u
MI16 Z net25 VSS VSS nch w=0.39u l=0.06u
MI8_1 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_2 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_0 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI21 net024 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHD2 I Z VDD VDDL VSS
MI15_0 VDD net25 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net25 Z VDD pch w=0.52u l=0.06u
MI5 VDD net25 net34 VDD pch w=0.15u l=0.06u
MI19 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI17 net25 net34 VDD VDD pch w=0.15u l=0.06u
MI6_0 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_1 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_2 net25 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z net25 VSS VSS nch w=0.39u l=0.06u
MI8_0 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_1 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z net25 VSS VSS nch w=0.39u l=0.06u
MI21 net024 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHD4 I Z VDD VDDL VSS
MI15_0 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD p0 Z VDD pch w=0.52u l=0.06u
MI5 VDD p0 net031 VDD pch w=0.15u l=0.06u
MI19 net49 I VDDL VDDL pch w=0.52u l=0.06u
MI17 p0 net031 VDD VDD pch w=0.15u l=0.06u
MI6_0 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_1 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_2 p0 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_3 Z p0 VSS VSS nch w=0.39u l=0.06u
MI8_0 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_1 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI21 net49 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHD8 I Z VDD VDDL VSS
MI15_0 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_4 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_5 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_6 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_7 VDD p0 Z VDD pch w=0.52u l=0.06u
MI5 VDD p0 net031 VDD pch w=0.15u l=0.06u
MI19 net49 I VDDL VDDL pch w=0.52u l=0.06u
MI17 p0 net031 VDD VDD pch w=0.15u l=0.06u
MI6_0 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_1 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_2 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_3 p0 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_3 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_4 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_5 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_6 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_7 Z p0 VSS VSS nch w=0.39u l=0.06u
MI8_0 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_1 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_2 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI21 net49 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFACD1 I NSLEEP Z VDD VDDL VSS
MI16 Z net031 vvss VSS nch w=0.39u l=0.06u
MI44 net024 I vvss VSS nch w=0.39u l=0.06u
MI43_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI43_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI43_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40_0 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_1 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_2 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_3 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI42_0 net031 I vvss VSS nch w=0.39u l=0.06u
MI42_1 net031 I vvss VSS nch w=0.39u l=0.06u
MI42_2 net031 I vvss VSS nch w=0.39u l=0.06u
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net031 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net031 net34 VDD pch w=0.15u l=0.06u
MI15 VDD net031 Z VDD pch w=0.52u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.15u l=0.06u
.ends
.subckt LVLLHFACD2 I NSLEEP Z VDD VDDL VSS
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net043 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net043 net34 VDD pch w=0.15u l=0.06u
MI15_0 VDD net043 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net043 Z VDD pch w=0.52u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.34u l=0.06u
MI16_0 Z net043 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net043 vvss VSS nch w=0.39u l=0.06u
MI45 net024 I vvss VSS nch w=0.39u l=0.06u
MI44_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI44_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI44_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40_0 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_1 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_2 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI40_3 vvss NSLEEP VSS VSS nch w=0.39u l=0.06u
MI43_0 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_1 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_2 net043 I vvss VSS nch w=0.39u l=0.06u
MI43_3 net043 I vvss VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFACD4 I NSLEEP Z VDD VDDL VSS
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net038 net34 VDD VDD pch w=0.15u l=0.06u
MI15_0 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD net038 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD net038 Z VDD pch w=0.52u l=0.06u
MI37 VDD net038 net34 VDD pch w=0.15u l=0.06u
MI41 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
MI45_0 net038 I vvss VSS nch w=0.39u l=0.06u
MI45_1 net038 I vvss VSS nch w=0.39u l=0.06u
MI45_2 net038 I vvss VSS nch w=0.39u l=0.06u
MI46_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI40 vvss NSLEEP VSS VSS nch w=3.11u l=0.06u
MI16_0 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_2 Z net038 vvss VSS nch w=0.39u l=0.06u
MI16_3 Z net038 vvss VSS nch w=0.39u l=0.06u
MI47 net024 I vvss VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFACD8 I NSLEEP Z VDD VDDL VSS
MI45_0 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_1 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_2 net087 I vvss VSS nch w=0.39u l=0.06u
MI45_3 net087 I vvss VSS nch w=0.39u l=0.06u
MI46_0 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_1 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI46_2 net34 net024 vvss VSS nch w=0.39u l=0.06u
MI16_0 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_1 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_2 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_3 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_4 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_5 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_6 Z net087 vvss VSS nch w=0.39u l=0.06u
MI16_7 Z net087 vvss VSS nch w=0.39u l=0.06u
MI40 vvss NSLEEP VSS VSS nch w=6.26u l=0.06u
MI47 net024 I vvss VSS nch w=0.39u l=0.06u
MI33 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI36 net087 net34 VDD VDD pch w=0.15u l=0.06u
MI37 VDD net087 net34 VDD pch w=0.15u l=0.06u
MI15_0 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_4 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_5 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_6 VDD net087 Z VDD pch w=0.52u l=0.06u
MI15_7 VDD net087 Z VDD pch w=0.52u l=0.06u
MI41_0 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
MI41_1 Z NSLEEP VDD VDD pch w=0.52u l=0.06u
.ends
.subckt LVLLHFAD1 I Z VDD VDDL VSS
MI15 VDD net25 Z VDD pch w=0.52u l=0.06u
MI5 VDD net25 net34 VDD pch w=0.15u l=0.06u
MI19 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI17 net25 net34 VDD VDD pch w=0.15u l=0.06u
MI6_0 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_1 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_2 net25 I VSS VSS nch w=0.39u l=0.06u
MI16 Z net25 VSS VSS nch w=0.39u l=0.06u
MI8_1 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_2 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_0 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI21 net024 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFAD2 I Z VDD VDDL VSS
MI15_0 VDD net25 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD net25 Z VDD pch w=0.52u l=0.06u
MI5 VDD net25 net34 VDD pch w=0.15u l=0.06u
MI19 net024 I VDDL VDDL pch w=0.52u l=0.06u
MI17 net25 net34 VDD VDD pch w=0.15u l=0.06u
MI6_0 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_1 net25 I VSS VSS nch w=0.39u l=0.06u
MI6_2 net25 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z net25 VSS VSS nch w=0.39u l=0.06u
MI8_0 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI8_1 net34 net024 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z net25 VSS VSS nch w=0.39u l=0.06u
MI21 net024 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFAD4 I Z VDD VDDL VSS
MI15_0 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD p0 Z VDD pch w=0.52u l=0.06u
MI5 VDD p0 net031 VDD pch w=0.15u l=0.06u
MI19 net49 I VDDL VDDL pch w=0.52u l=0.06u
MI17 p0 net031 VDD VDD pch w=0.15u l=0.06u
MI6_0 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_1 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_2 p0 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_3 Z p0 VSS VSS nch w=0.39u l=0.06u
MI8_0 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_1 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI21 net49 I VSS VSS nch w=0.39u l=0.06u
.ends
.subckt LVLLHFAD8 I Z VDD VDDL VSS
MI15_0 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_1 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_2 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_3 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_4 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_5 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_6 VDD p0 Z VDD pch w=0.52u l=0.06u
MI15_7 VDD p0 Z VDD pch w=0.52u l=0.06u
MI5 VDD p0 net031 VDD pch w=0.15u l=0.06u
MI19 net49 I VDDL VDDL pch w=0.52u l=0.06u
MI17 p0 net031 VDD VDD pch w=0.15u l=0.06u
MI6_0 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_1 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_2 p0 I VSS VSS nch w=0.39u l=0.06u
MI6_3 p0 I VSS VSS nch w=0.39u l=0.06u
MI16_0 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_1 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_2 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_3 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_4 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_5 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_6 Z p0 VSS VSS nch w=0.39u l=0.06u
MI16_7 Z p0 VSS VSS nch w=0.39u l=0.06u
MI8_0 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_1 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI8_2 net031 net49 VSS VSS nch w=0.39u l=0.06u
MI21 net49 I VSS VSS nch w=0.39u l=0.06u
.ends
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        