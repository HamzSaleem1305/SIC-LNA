magic
tech sky130A
magscale 1 2
timestamp 1666417074
<< pwell >>
rect 6500 -670 7960 440
rect 3130 -2610 7960 -670
rect 6500 -5040 7960 -2610
<< ndiff >>
rect 6192 -2118 6286 -2102
<< poly >>
rect 5030 -870 5640 -800
rect 6190 -1360 6420 -1290
rect 5010 -2270 5660 -2200
rect 6170 -2270 6430 -2200
<< locali >>
rect 7170 400 7785 435
rect 7170 250 7520 400
rect 7660 250 7785 400
rect 7170 225 7785 250
rect 4870 -2170 5020 -2040
rect 7170 -2080 7380 225
rect 7170 -2170 7190 -2080
rect 7360 -2170 7380 -2080
rect 6900 -2910 7060 -2560
rect 7170 -4060 7380 -2170
rect 7170 -5200 7390 -4060
rect 7090 -5280 7390 -5200
<< viali >>
rect 7520 250 7660 400
rect 7190 -2170 7360 -2080
<< metal1 >>
rect 7500 400 7680 430
rect 7500 250 7520 400
rect 7660 250 7680 400
rect 7500 30 7680 250
rect 6930 -430 7280 10
rect 7540 -270 7630 30
rect 5030 -790 5640 -770
rect 5030 -850 5070 -790
rect 5610 -850 5640 -790
rect 5030 -860 5640 -850
rect 5050 -910 5130 -900
rect 5050 -1020 5060 -910
rect 5120 -1020 5130 -910
rect 5050 -1030 5130 -1020
rect 5240 -910 5320 -900
rect 5240 -1020 5250 -910
rect 5310 -1020 5320 -910
rect 5240 -1030 5320 -1020
rect 5440 -910 5520 -900
rect 5440 -1020 5450 -910
rect 5510 -1020 5520 -910
rect 5440 -1030 5520 -1020
rect 5630 -910 5710 -900
rect 5630 -1020 5640 -910
rect 5700 -1020 5710 -910
rect 5630 -1030 5710 -1020
rect 6270 -1350 6330 -1290
rect 6210 -1390 6290 -1380
rect 6210 -1500 6220 -1390
rect 6280 -1500 6290 -1390
rect 6210 -1510 6290 -1500
rect 6400 -1390 6480 -1380
rect 6400 -1500 6410 -1390
rect 6470 -1500 6480 -1390
rect 6400 -1510 6480 -1500
rect 4960 -2050 5040 -2040
rect 4960 -2160 4970 -2050
rect 5030 -2160 5040 -2050
rect 4960 -2170 5040 -2160
rect 5150 -2050 5230 -2040
rect 5150 -2160 5160 -2050
rect 5220 -2160 5230 -2050
rect 5150 -2170 5230 -2160
rect 5340 -2050 5420 -2040
rect 5340 -2160 5350 -2050
rect 5410 -2160 5420 -2050
rect 5340 -2170 5420 -2160
rect 5530 -2050 5610 -2040
rect 5530 -2160 5540 -2050
rect 5600 -2160 5610 -2050
rect 5530 -2170 5610 -2160
rect 6110 -2060 6190 -2050
rect 6110 -2170 6120 -2060
rect 6180 -2170 6190 -2060
rect 6110 -2180 6190 -2170
rect 6310 -2060 6390 -2050
rect 6310 -2170 6320 -2060
rect 6380 -2170 6390 -2060
rect 6310 -2180 6390 -2170
rect 7170 -2080 7380 -2060
rect 7170 -2170 7190 -2080
rect 7360 -2170 7380 -2080
rect 7170 -2180 7380 -2170
rect 5010 -2280 5660 -2210
rect 6170 -2220 6760 -2210
rect 6170 -2270 6650 -2220
rect 5290 -2360 5410 -2280
rect 6640 -2310 6650 -2270
rect 6750 -2310 6760 -2220
rect 6640 -2320 6760 -2310
rect 5290 -2480 7010 -2360
rect 6930 -3300 7030 -2990
rect 6930 -3400 6940 -3300
rect 7020 -3400 7030 -3300
rect 6930 -3410 7030 -3400
rect 7480 -3300 7680 -3280
rect 5930 -3730 7130 -3470
rect 7480 -3600 7500 -3300
rect 7660 -3600 7680 -3300
rect 7480 -3620 7680 -3600
rect 6870 -3810 7130 -3730
rect 6870 -4040 6910 -3810
rect 7100 -4040 7130 -3810
rect 6870 -4070 7130 -4040
<< via1 >>
rect 5070 -850 5610 -790
rect 5060 -1020 5120 -910
rect 5250 -1020 5310 -910
rect 5450 -1020 5510 -910
rect 5640 -1020 5700 -910
rect 6220 -1500 6280 -1390
rect 6410 -1500 6470 -1390
rect 4970 -2160 5030 -2050
rect 5160 -2160 5220 -2050
rect 5350 -2160 5410 -2050
rect 5540 -2160 5600 -2050
rect 6120 -2170 6180 -2060
rect 6320 -2170 6380 -2060
rect 7190 -2170 7360 -2080
rect 6650 -2310 6750 -2220
rect 6940 -3400 7020 -3300
rect 7500 -3600 7660 -3300
rect 6910 -4040 7100 -3810
<< metal2 >>
rect 4690 -790 5640 -770
rect 4690 -850 5070 -790
rect 5610 -850 5640 -790
rect 4690 -870 5640 -850
rect 4700 -1320 4800 -870
rect 5050 -910 5895 -900
rect 5050 -1020 5060 -910
rect 5120 -1020 5250 -910
rect 5310 -1020 5450 -910
rect 5510 -1020 5640 -910
rect 5700 -1020 5895 -910
rect 5050 -1030 5895 -1020
rect 3160 -1420 4800 -1320
rect 5765 -1375 5895 -1030
rect 5765 -1380 6325 -1375
rect 5765 -1390 6480 -1380
rect 2790 -4240 3090 -4210
rect 2790 -4480 2810 -4240
rect 3060 -4260 3090 -4240
rect 3160 -4260 3260 -1420
rect 5765 -1500 6220 -1390
rect 6280 -1500 6410 -1390
rect 6470 -1500 6480 -1390
rect 5765 -1505 6325 -1500
rect 6210 -1510 6290 -1505
rect 6400 -1510 6480 -1500
rect 4960 -2050 5610 -2040
rect 4960 -2160 4970 -2050
rect 5030 -2160 5160 -2050
rect 5220 -2160 5350 -2050
rect 5410 -2160 5540 -2050
rect 5600 -2160 5610 -2050
rect 4960 -2170 5610 -2160
rect 6110 -2060 6190 -2050
rect 6310 -2060 6390 -2050
rect 6110 -2170 6120 -2060
rect 6180 -2170 6320 -2060
rect 6380 -2080 7380 -2060
rect 6380 -2170 7190 -2080
rect 7360 -2170 7380 -2080
rect 6110 -2180 7380 -2170
rect 6640 -2220 6770 -2210
rect 6640 -2310 6650 -2220
rect 6750 -2310 6770 -2220
rect 6640 -2320 6770 -2310
rect 6650 -3290 6770 -2320
rect 8350 -2270 8740 -2230
rect 8350 -2355 8380 -2270
rect 7875 -2645 8380 -2355
rect 7480 -3290 7680 -3280
rect 6650 -3300 7680 -3290
rect 6650 -3400 6940 -3300
rect 7020 -3400 7500 -3300
rect 6650 -3410 7500 -3400
rect 7480 -3600 7500 -3410
rect 7660 -3600 7680 -3300
rect 7480 -3620 7680 -3600
rect 7875 -3770 8165 -2645
rect 8350 -2730 8380 -2645
rect 8710 -2355 8740 -2270
rect 8710 -2645 8785 -2355
rect 8710 -2730 8740 -2645
rect 8350 -2760 8740 -2730
rect 6870 -3774 7380 -3770
rect 7420 -3774 8170 -3770
rect 6870 -3810 8170 -3774
rect 6870 -4040 6910 -3810
rect 7100 -4040 8170 -3810
rect 6870 -4054 8170 -4040
rect 6870 -4060 7380 -4054
rect 7420 -4060 8170 -4054
rect 3060 -4360 3260 -4260
rect 3060 -4480 3090 -4360
rect 2790 -4510 3090 -4480
rect 3010 -4786 4596 -4626
rect 2640 -5230 2920 -5200
rect 2640 -5550 2660 -5230
rect 2900 -5340 2920 -5230
rect 3010 -5340 3170 -4786
rect 2900 -5500 3170 -5340
rect 2900 -5550 2920 -5500
rect 2640 -5570 2920 -5550
<< via2 >>
rect 2810 -4480 3060 -4240
rect 7500 -3600 7660 -3300
rect 8380 -2730 8710 -2270
rect 2660 -5550 2900 -5230
<< metal3 >>
rect 8350 -2270 8740 -2230
rect 8350 -2730 8380 -2270
rect 8710 -2730 8740 -2270
rect 8350 -2760 8740 -2730
rect 7480 -3300 7680 -3280
rect 7480 -3600 7500 -3300
rect 7660 -3600 7680 -3300
rect 7480 -3620 7680 -3600
rect 2790 -4240 3090 -4210
rect 2790 -4480 2810 -4240
rect 3060 -4480 3090 -4240
rect 2790 -4510 3090 -4480
rect 2640 -5230 2920 -5200
rect 2640 -5550 2660 -5230
rect 2900 -5550 2920 -5230
rect 2640 -5570 2920 -5550
<< via3 >>
rect 8380 -2730 8710 -2270
rect 7500 -3600 7660 -3300
rect 2810 -4480 3060 -4240
rect 2660 -5550 2900 -5230
<< metal4 >>
rect 8350 -2270 8740 -2230
rect 8350 -2730 8380 -2270
rect 8710 -2730 8740 -2270
rect 8350 -2760 8740 -2730
rect 7480 -3300 9390 -3280
rect 7480 -3600 7500 -3300
rect 7660 -3600 9390 -3300
rect 7480 -3620 9390 -3600
rect 2210 -4240 3090 -4210
rect 2210 -4480 2810 -4240
rect 3060 -4480 3090 -4240
rect 2210 -4510 3090 -4480
rect 2640 -5230 2920 -5200
rect 2640 -5550 2660 -5230
rect 2900 -5550 2920 -5230
rect 2640 -5570 2920 -5550
<< via4 >>
rect 8380 -2730 8710 -2270
rect 2660 -5550 2900 -5230
<< metal5 >>
rect 8350 -2270 9410 -2230
rect 8350 -2730 8380 -2270
rect 8710 -2730 9410 -2270
rect 8350 -2760 9410 -2730
rect 2020 -5230 2950 -5180
rect 2020 -5550 2660 -5230
rect 2900 -5550 2950 -5230
rect 2020 -5590 2950 -5550
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC7
timestamp 1666381508
transform 0 1 12111 -1 0 -237
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC8
timestamp 1666381508
transform 0 -1 -759 1 0 -7559
box -3351 -3101 3373 3101
use sky130_fd_pr__nfet_01v8_lvt_2SWTDU  XM17
timestamp 1666381508
transform 1 0 5333 0 1 -1537
box -503 -853 503 853
use sky130_fd_pr__nfet_01v8_lvt_95PS5T  XM18
timestamp 1666381508
transform 1 0 6301 0 1 -1780
box -311 -610 311 610
use sky130_fd_pr__res_high_po_0p35_MTHP3S  XR11
timestamp 1666381508
transform 1 0 7581 0 1 -1902
box -201 -2098 201 2098
use sky130_fd_pr__res_high_po_0p35_M3EX2E  XR12
timestamp 1666381508
transform 1 0 6971 0 1 -1222
box -201 -1398 201 1398
use partition2  partition2_0
timestamp 1666417074
transform 1 0 -8194 0 1 -11626
box 11324 526 23405 10182
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1666383890
transform 1 0 6983 0 1 -3027
box -183 -183 183 183
<< labels >>
flabel metal1 7200 -220 7200 -220 0 FreeSans 800 0 0 0 VB0_9
flabel metal2 5840 -1150 5840 -1150 0 FreeSans 800 0 0 0 Vo2
flabel locali 7378 332 7378 332 0 FreeSans 1600 0 0 0 VDD
<< end >>
