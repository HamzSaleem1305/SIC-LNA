magic
tech sky130A
magscale 1 2
timestamp 1666417074
<< error_p >>
rect -29 1081 29 1087
rect -29 1047 -17 1081
rect -29 1041 29 1047
rect -125 -1047 -67 -1041
rect 67 -1047 125 -1041
rect -125 -1081 -113 -1047
rect 67 -1081 79 -1047
rect -125 -1087 -67 -1081
rect 67 -1087 125 -1081
<< nwell >>
rect -311 -1219 311 1219
<< pmos >>
rect -111 -1000 -81 1000
rect -15 -1000 15 1000
rect 81 -1000 111 1000
<< pdiff >>
rect -173 988 -111 1000
rect -173 -988 -161 988
rect -127 -988 -111 988
rect -173 -1000 -111 -988
rect -81 988 -15 1000
rect -81 -988 -65 988
rect -31 -988 -15 988
rect -81 -1000 -15 -988
rect 15 988 81 1000
rect 15 -988 31 988
rect 65 -988 81 988
rect 15 -1000 81 -988
rect 111 988 173 1000
rect 111 -988 127 988
rect 161 -988 173 988
rect 111 -1000 173 -988
<< pdiffc >>
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
<< nsubdiff >>
rect -275 1149 -179 1183
rect 179 1149 275 1183
rect -275 1087 -241 1149
rect 241 1087 275 1149
rect -275 -1149 -241 -1087
rect 241 -1149 275 -1087
rect -275 -1183 -179 -1149
rect 179 -1183 275 -1149
<< nsubdiffcont >>
rect -179 1149 179 1183
rect -275 -1087 -241 1087
rect 241 -1087 275 1087
rect -179 -1183 179 -1149
<< poly >>
rect -33 1081 33 1097
rect -33 1047 -17 1081
rect 17 1047 33 1081
rect -33 1031 33 1047
rect -111 1000 -81 1026
rect -15 1000 15 1031
rect 81 1000 111 1026
rect -111 -1031 -81 -1000
rect -15 -1026 15 -1000
rect 81 -1031 111 -1000
rect -129 -1047 -63 -1031
rect -129 -1081 -113 -1047
rect -79 -1081 -63 -1047
rect -129 -1097 -63 -1081
rect 63 -1047 129 -1031
rect 63 -1081 79 -1047
rect 113 -1081 129 -1047
rect 63 -1097 129 -1081
<< polycont >>
rect -17 1047 17 1081
rect -113 -1081 -79 -1047
rect 79 -1081 113 -1047
<< locali >>
rect -275 1149 -179 1183
rect 179 1149 275 1183
rect -275 1087 -241 1149
rect 241 1087 275 1149
rect -33 1047 -17 1081
rect 17 1047 33 1081
rect -161 988 -127 1004
rect -161 -1004 -127 -988
rect -65 988 -31 1004
rect -65 -1004 -31 -988
rect 31 988 65 1004
rect 31 -1004 65 -988
rect 127 988 161 1004
rect 127 -1004 161 -988
rect -129 -1081 -113 -1047
rect -79 -1081 -63 -1047
rect 63 -1081 79 -1047
rect 113 -1081 129 -1047
rect -275 -1149 -241 -1087
rect 241 -1149 275 -1087
rect -275 -1183 -179 -1149
rect 179 -1183 275 -1149
<< viali >>
rect -17 1047 17 1081
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
rect -113 -1081 -79 -1047
rect 79 -1081 113 -1047
<< metal1 >>
rect -29 1081 29 1087
rect -29 1047 -17 1081
rect 17 1047 29 1081
rect -29 1041 29 1047
rect -167 988 -121 1000
rect -167 -988 -161 988
rect -127 -988 -121 988
rect -167 -1000 -121 -988
rect -71 988 -25 1000
rect -71 -988 -65 988
rect -31 -988 -25 988
rect -71 -1000 -25 -988
rect 25 988 71 1000
rect 25 -988 31 988
rect 65 -988 71 988
rect 25 -1000 71 -988
rect 121 988 167 1000
rect 121 -988 127 988
rect 161 -988 167 988
rect 121 -1000 167 -988
rect -125 -1047 -67 -1041
rect -125 -1081 -113 -1047
rect -79 -1081 -67 -1047
rect -125 -1087 -67 -1081
rect 67 -1047 125 -1041
rect 67 -1081 79 -1047
rect 113 -1081 125 -1047
rect 67 -1087 125 -1081
<< properties >>
string FIXED_BBOX -258 -1166 258 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
