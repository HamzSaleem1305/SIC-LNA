magic
tech sky130A
magscale 1 2
timestamp 1666374491
<< pwell >>
rect -235 -667 235 667
<< psubdiff >>
rect -199 597 -103 631
rect 103 597 199 631
rect -199 535 -165 597
rect 165 535 199 597
rect -199 -597 -165 -535
rect 165 -597 199 -535
rect -199 -631 -103 -597
rect 103 -631 199 -597
<< psubdiffcont >>
rect -103 597 103 631
rect -199 -535 -165 535
rect 165 -535 199 535
rect -103 -631 103 -597
<< xpolycontact >>
rect -69 69 69 501
rect -69 -501 69 -69
<< ppolyres >>
rect -69 -69 69 69
<< locali >>
rect -199 597 -103 631
rect 103 597 199 631
rect -199 535 -165 597
rect 165 535 199 597
rect -199 -597 -165 -535
rect 165 -597 199 -535
rect -199 -631 -103 -597
rect 103 -631 199 -597
<< viali >>
rect -53 86 53 483
rect -53 -483 53 -86
<< metal1 >>
rect -59 483 59 495
rect -59 86 -53 483
rect 53 86 59 483
rect -59 74 59 86
rect -59 -86 59 -74
rect -59 -483 -53 -86
rect 53 -483 59 -86
rect -59 -495 59 -483
<< res0p69 >>
rect -71 -71 71 71
<< properties >>
string FIXED_BBOX -182 -614 182 614
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.69 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 375.417 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
