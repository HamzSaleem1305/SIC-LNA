magic
tech sky130A
magscale 1 2
timestamp 1666374491
<< pwell >>
rect -1586 -667 1586 667
<< psubdiff >>
rect -1550 597 -1454 631
rect 1454 597 1550 631
rect -1550 535 -1516 597
rect 1516 535 1550 597
rect -1550 -597 -1516 -535
rect 1516 -597 1550 -535
rect -1550 -631 -1454 -597
rect 1454 -631 1550 -597
<< psubdiffcont >>
rect -1454 597 1454 631
rect -1550 -535 -1516 535
rect 1516 -535 1550 535
rect -1454 -631 1454 -597
<< xpolycontact >>
rect -1420 69 -1282 501
rect -1420 -501 -1282 -69
rect -1034 69 -896 501
rect -1034 -501 -896 -69
rect -648 69 -510 501
rect -648 -501 -510 -69
rect -262 69 -124 501
rect -262 -501 -124 -69
rect 124 69 262 501
rect 124 -501 262 -69
rect 510 69 648 501
rect 510 -501 648 -69
rect 896 69 1034 501
rect 896 -501 1034 -69
rect 1282 69 1420 501
rect 1282 -501 1420 -69
<< ppolyres >>
rect -1420 -69 -1282 69
rect -1034 -69 -896 69
rect -648 -69 -510 69
rect -262 -69 -124 69
rect 124 -69 262 69
rect 510 -69 648 69
rect 896 -69 1034 69
rect 1282 -69 1420 69
<< locali >>
rect -1550 597 -1454 631
rect 1454 597 1550 631
rect -1550 535 -1516 597
rect 1516 535 1550 597
rect -1550 -597 -1516 -535
rect 1516 -597 1550 -535
rect -1550 -631 -1454 -597
rect 1454 -631 1550 -597
<< viali >>
rect -1404 86 -1298 483
rect -1018 86 -912 483
rect -632 86 -526 483
rect -246 86 -140 483
rect 140 86 246 483
rect 526 86 632 483
rect 912 86 1018 483
rect 1298 86 1404 483
rect -1404 -483 -1298 -86
rect -1018 -483 -912 -86
rect -632 -483 -526 -86
rect -246 -483 -140 -86
rect 140 -483 246 -86
rect 526 -483 632 -86
rect 912 -483 1018 -86
rect 1298 -483 1404 -86
<< metal1 >>
rect -1410 483 -1292 495
rect -1410 86 -1404 483
rect -1298 86 -1292 483
rect -1410 74 -1292 86
rect -1024 483 -906 495
rect -1024 86 -1018 483
rect -912 86 -906 483
rect -1024 74 -906 86
rect -638 483 -520 495
rect -638 86 -632 483
rect -526 86 -520 483
rect -638 74 -520 86
rect -252 483 -134 495
rect -252 86 -246 483
rect -140 86 -134 483
rect -252 74 -134 86
rect 134 483 252 495
rect 134 86 140 483
rect 246 86 252 483
rect 134 74 252 86
rect 520 483 638 495
rect 520 86 526 483
rect 632 86 638 483
rect 520 74 638 86
rect 906 483 1024 495
rect 906 86 912 483
rect 1018 86 1024 483
rect 906 74 1024 86
rect 1292 483 1410 495
rect 1292 86 1298 483
rect 1404 86 1410 483
rect 1292 74 1410 86
rect -1410 -86 -1292 -74
rect -1410 -483 -1404 -86
rect -1298 -483 -1292 -86
rect -1410 -495 -1292 -483
rect -1024 -86 -906 -74
rect -1024 -483 -1018 -86
rect -912 -483 -906 -86
rect -1024 -495 -906 -483
rect -638 -86 -520 -74
rect -638 -483 -632 -86
rect -526 -483 -520 -86
rect -638 -495 -520 -483
rect -252 -86 -134 -74
rect -252 -483 -246 -86
rect -140 -483 -134 -86
rect -252 -495 -134 -483
rect 134 -86 252 -74
rect 134 -483 140 -86
rect 246 -483 252 -86
rect 134 -495 252 -483
rect 520 -86 638 -74
rect 520 -483 526 -86
rect 632 -483 638 -86
rect 520 -495 638 -483
rect 906 -86 1024 -74
rect 906 -483 912 -86
rect 1018 -483 1024 -86
rect 906 -495 1024 -483
rect 1292 -86 1410 -74
rect 1292 -483 1298 -86
rect 1404 -483 1410 -86
rect 1292 -495 1410 -483
<< res0p69 >>
rect -1422 -71 -1280 71
rect -1036 -71 -894 71
rect -650 -71 -508 71
rect -264 -71 -122 71
rect 122 -71 264 71
rect 508 -71 650 71
rect 894 -71 1036 71
rect 1280 -71 1422 71
<< properties >>
string FIXED_BBOX -1533 -614 1533 614
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.69 m 1 nx 8 wmin 0.690 lmin 0.50 rho 319.8 val 375.417 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
