magic
tech sky130A
magscale 1 2
timestamp 1666476701
<< nwell >>
rect 15680 20970 16302 23408
rect 16942 13724 17564 16162
<< pwell >>
rect 12944 24782 15584 24787
rect 16341 24782 17808 24794
rect 12880 24380 17808 24782
rect 12944 24102 15584 24380
rect 12910 23700 15584 24102
rect 12944 23390 15584 23700
rect 12944 22943 15600 23390
rect 12980 20670 15600 22943
rect 16341 21780 17808 24380
rect 16341 21778 17810 21780
rect 16350 20670 17810 21778
rect 12980 18730 17810 20670
rect 12986 16300 17810 18730
rect 12986 13699 16476 16300
rect 12984 10534 17949 13699
<< pmos >>
rect 15880 21189 15910 23189
rect 15976 21189 16006 23189
rect 16072 21189 16102 23189
rect 17142 13943 17172 15943
rect 17238 13943 17268 15943
rect 17334 13943 17364 15943
<< nmoslvt >>
rect 14020 21150 14050 23150
rect 14116 21150 14146 23150
rect 14212 21150 14242 23150
rect 14308 21150 14338 23150
rect 14404 21150 14434 23150
rect 14500 21150 14530 23150
rect 14596 21150 14626 23150
rect 14692 21150 14722 23150
rect 16712 22040 16742 24040
rect 16808 22040 16838 24040
rect 16904 22040 16934 24040
rect 17000 22040 17030 24040
rect 17096 22040 17126 24040
rect 17192 22040 17222 24040
rect 17288 22040 17318 24040
rect 17384 22040 17414 24040
rect 17480 22040 17510 24040
rect 17576 22040 17606 24040
rect 14880 19160 14910 20446
rect 14976 19160 15006 20446
rect 15072 19160 15102 20446
rect 15168 19160 15198 20446
rect 15264 19160 15294 20446
rect 15360 19160 15390 20446
rect 15456 19160 15486 20446
rect 16040 19160 16070 19960
rect 16136 19160 16166 19960
rect 16232 19160 16262 19960
rect 15062 16934 15092 18494
rect 15472 16934 15502 18494
rect 13618 13904 13648 15464
rect 14472 13904 14502 15904
rect 14568 13904 14598 15904
rect 14664 13904 14694 15904
rect 14760 13904 14790 15904
rect 14856 13904 14886 15904
rect 14952 13904 14982 15904
rect 15048 13904 15078 15904
rect 15144 13904 15174 15904
rect 13480 11070 13510 13070
rect 13568 11070 13598 13070
rect 13656 11070 13686 13070
rect 13744 11070 13774 13070
rect 13832 11070 13862 13070
rect 13920 11070 13950 13070
rect 14008 11070 14038 13070
rect 14096 11070 14126 13070
rect 14184 11070 14214 13070
rect 14272 11070 14302 13070
rect 14360 11070 14390 13070
rect 14448 11070 14478 13070
rect 14536 11070 14566 13070
rect 14624 11070 14654 13070
rect 14712 11070 14742 13070
rect 14800 11070 14830 13070
rect 14888 11070 14918 13070
rect 14976 11070 15006 13070
rect 15064 11070 15094 13070
rect 15152 11070 15182 13070
rect 15240 11070 15270 13070
rect 15328 11070 15358 13070
rect 15416 11070 15446 13070
rect 15504 11070 15534 13070
rect 15592 11070 15622 13070
rect 15680 11070 15710 13070
rect 15768 11070 15798 13070
rect 15856 11070 15886 13070
rect 15944 11070 15974 13070
rect 16032 11070 16062 13070
rect 16120 11070 16150 13070
rect 16208 11070 16238 13070
rect 16296 11070 16326 13070
rect 16384 11070 16414 13070
rect 16472 11070 16502 13070
rect 16560 11070 16590 13070
rect 16648 11070 16678 13070
rect 16736 11070 16766 13070
rect 16824 11070 16854 13070
rect 16912 11070 16942 13070
rect 17000 11070 17030 13070
rect 17088 11070 17118 13070
rect 17176 11070 17206 13070
rect 17264 11070 17294 13070
rect 17352 11070 17382 13070
rect 17440 11070 17470 13070
<< ndiff >>
rect 13958 23138 14020 23150
rect 13958 21162 13970 23138
rect 14004 21162 14020 23138
rect 13958 21150 14020 21162
rect 14050 23138 14116 23150
rect 14050 21162 14066 23138
rect 14100 21162 14116 23138
rect 14050 21150 14116 21162
rect 14146 23138 14212 23150
rect 14146 21162 14162 23138
rect 14196 21162 14212 23138
rect 14146 21150 14212 21162
rect 14242 23138 14308 23150
rect 14242 21162 14258 23138
rect 14292 21162 14308 23138
rect 14242 21150 14308 21162
rect 14338 23138 14404 23150
rect 14338 21162 14354 23138
rect 14388 21162 14404 23138
rect 14338 21150 14404 21162
rect 14434 23138 14500 23150
rect 14434 21162 14450 23138
rect 14484 21162 14500 23138
rect 14434 21150 14500 21162
rect 14530 23138 14596 23150
rect 14530 21162 14546 23138
rect 14580 21162 14596 23138
rect 14530 21150 14596 21162
rect 14626 23138 14692 23150
rect 14626 21162 14642 23138
rect 14676 21162 14692 23138
rect 14626 21150 14692 21162
rect 14722 23138 14784 23150
rect 14722 21162 14738 23138
rect 14772 21162 14784 23138
rect 14722 21150 14784 21162
rect 16650 24028 16712 24040
rect 16650 22052 16662 24028
rect 16696 22052 16712 24028
rect 16650 22040 16712 22052
rect 16742 24028 16808 24040
rect 16742 22052 16758 24028
rect 16792 22052 16808 24028
rect 16742 22040 16808 22052
rect 16838 24028 16904 24040
rect 16838 22052 16854 24028
rect 16888 22052 16904 24028
rect 16838 22040 16904 22052
rect 16934 24028 17000 24040
rect 16934 22052 16950 24028
rect 16984 22052 17000 24028
rect 16934 22040 17000 22052
rect 17030 24028 17096 24040
rect 17030 22052 17046 24028
rect 17080 22052 17096 24028
rect 17030 22040 17096 22052
rect 17126 24028 17192 24040
rect 17126 22052 17142 24028
rect 17176 22052 17192 24028
rect 17126 22040 17192 22052
rect 17222 24028 17288 24040
rect 17222 22052 17238 24028
rect 17272 22052 17288 24028
rect 17222 22040 17288 22052
rect 17318 24028 17384 24040
rect 17318 22052 17334 24028
rect 17368 22052 17384 24028
rect 17318 22040 17384 22052
rect 17414 24028 17480 24040
rect 17414 22052 17430 24028
rect 17464 22052 17480 24028
rect 17414 22040 17480 22052
rect 17510 24028 17576 24040
rect 17510 22052 17526 24028
rect 17560 22052 17576 24028
rect 17510 22040 17576 22052
rect 17606 24028 17668 24040
rect 17606 22052 17622 24028
rect 17656 22052 17668 24028
rect 17606 22040 17668 22052
rect 14818 20434 14880 20446
rect 14818 19172 14830 20434
rect 14864 19172 14880 20434
rect 14818 19160 14880 19172
rect 14910 20434 14976 20446
rect 14910 19172 14926 20434
rect 14960 19172 14976 20434
rect 14910 19160 14976 19172
rect 15006 20434 15072 20446
rect 15006 19172 15022 20434
rect 15056 19172 15072 20434
rect 15006 19160 15072 19172
rect 15102 20434 15168 20446
rect 15102 19172 15118 20434
rect 15152 19172 15168 20434
rect 15102 19160 15168 19172
rect 15198 20434 15264 20446
rect 15198 19172 15214 20434
rect 15248 19172 15264 20434
rect 15198 19160 15264 19172
rect 15294 20434 15360 20446
rect 15294 19172 15310 20434
rect 15344 19172 15360 20434
rect 15294 19160 15360 19172
rect 15390 20434 15456 20446
rect 15390 19172 15406 20434
rect 15440 19172 15456 20434
rect 15390 19160 15456 19172
rect 15486 20434 15548 20446
rect 15486 19172 15502 20434
rect 15536 19172 15548 20434
rect 15486 19160 15548 19172
rect 15978 19948 16040 19960
rect 15978 19172 15990 19948
rect 16024 19172 16040 19948
rect 15978 19160 16040 19172
rect 16070 19948 16136 19960
rect 16070 19172 16086 19948
rect 16120 19172 16136 19948
rect 16070 19160 16136 19172
rect 16166 19948 16232 19960
rect 16166 19172 16182 19948
rect 16216 19172 16232 19948
rect 16166 19160 16232 19172
rect 16262 19948 16324 19960
rect 16262 19172 16278 19948
rect 16312 19172 16324 19948
rect 16262 19160 16324 19172
rect 15004 18482 15062 18494
rect 15004 16946 15016 18482
rect 15050 16946 15062 18482
rect 15004 16934 15062 16946
rect 15092 18482 15150 18494
rect 15092 16946 15104 18482
rect 15138 16946 15150 18482
rect 15092 16934 15150 16946
rect 15414 18482 15472 18494
rect 15414 16946 15426 18482
rect 15460 16946 15472 18482
rect 15414 16934 15472 16946
rect 15502 18482 15560 18494
rect 15502 16946 15514 18482
rect 15548 16946 15560 18482
rect 15502 16934 15560 16946
rect 13560 15452 13618 15464
rect 13560 13916 13572 15452
rect 13606 13916 13618 15452
rect 13560 13904 13618 13916
rect 13648 15452 13706 15464
rect 13648 13916 13660 15452
rect 13694 13916 13706 15452
rect 13648 13904 13706 13916
rect 14410 15892 14472 15904
rect 14410 13916 14422 15892
rect 14456 13916 14472 15892
rect 14410 13904 14472 13916
rect 14502 15892 14568 15904
rect 14502 13916 14518 15892
rect 14552 13916 14568 15892
rect 14502 13904 14568 13916
rect 14598 15892 14664 15904
rect 14598 13916 14614 15892
rect 14648 13916 14664 15892
rect 14598 13904 14664 13916
rect 14694 15892 14760 15904
rect 14694 13916 14710 15892
rect 14744 13916 14760 15892
rect 14694 13904 14760 13916
rect 14790 15892 14856 15904
rect 14790 13916 14806 15892
rect 14840 13916 14856 15892
rect 14790 13904 14856 13916
rect 14886 15892 14952 15904
rect 14886 13916 14902 15892
rect 14936 13916 14952 15892
rect 14886 13904 14952 13916
rect 14982 15892 15048 15904
rect 14982 13916 14998 15892
rect 15032 13916 15048 15892
rect 14982 13904 15048 13916
rect 15078 15892 15144 15904
rect 15078 13916 15094 15892
rect 15128 13916 15144 15892
rect 15078 13904 15144 13916
rect 15174 15892 15236 15904
rect 15174 13916 15190 15892
rect 15224 13916 15236 15892
rect 15174 13904 15236 13916
rect 13422 13058 13480 13070
rect 13422 11082 13434 13058
rect 13468 11082 13480 13058
rect 13422 11070 13480 11082
rect 13510 13058 13568 13070
rect 13510 11082 13522 13058
rect 13556 11082 13568 13058
rect 13510 11070 13568 11082
rect 13598 13058 13656 13070
rect 13598 11082 13610 13058
rect 13644 11082 13656 13058
rect 13598 11070 13656 11082
rect 13686 13058 13744 13070
rect 13686 11082 13698 13058
rect 13732 11082 13744 13058
rect 13686 11070 13744 11082
rect 13774 13058 13832 13070
rect 13774 11082 13786 13058
rect 13820 11082 13832 13058
rect 13774 11070 13832 11082
rect 13862 13058 13920 13070
rect 13862 11082 13874 13058
rect 13908 11082 13920 13058
rect 13862 11070 13920 11082
rect 13950 13058 14008 13070
rect 13950 11082 13962 13058
rect 13996 11082 14008 13058
rect 13950 11070 14008 11082
rect 14038 13058 14096 13070
rect 14038 11082 14050 13058
rect 14084 11082 14096 13058
rect 14038 11070 14096 11082
rect 14126 13058 14184 13070
rect 14126 11082 14138 13058
rect 14172 11082 14184 13058
rect 14126 11070 14184 11082
rect 14214 13058 14272 13070
rect 14214 11082 14226 13058
rect 14260 11082 14272 13058
rect 14214 11070 14272 11082
rect 14302 13058 14360 13070
rect 14302 11082 14314 13058
rect 14348 11082 14360 13058
rect 14302 11070 14360 11082
rect 14390 13058 14448 13070
rect 14390 11082 14402 13058
rect 14436 11082 14448 13058
rect 14390 11070 14448 11082
rect 14478 13058 14536 13070
rect 14478 11082 14490 13058
rect 14524 11082 14536 13058
rect 14478 11070 14536 11082
rect 14566 13058 14624 13070
rect 14566 11082 14578 13058
rect 14612 11082 14624 13058
rect 14566 11070 14624 11082
rect 14654 13058 14712 13070
rect 14654 11082 14666 13058
rect 14700 11082 14712 13058
rect 14654 11070 14712 11082
rect 14742 13058 14800 13070
rect 14742 11082 14754 13058
rect 14788 11082 14800 13058
rect 14742 11070 14800 11082
rect 14830 13058 14888 13070
rect 14830 11082 14842 13058
rect 14876 11082 14888 13058
rect 14830 11070 14888 11082
rect 14918 13058 14976 13070
rect 14918 11082 14930 13058
rect 14964 11082 14976 13058
rect 14918 11070 14976 11082
rect 15006 13058 15064 13070
rect 15006 11082 15018 13058
rect 15052 11082 15064 13058
rect 15006 11070 15064 11082
rect 15094 13058 15152 13070
rect 15094 11082 15106 13058
rect 15140 11082 15152 13058
rect 15094 11070 15152 11082
rect 15182 13058 15240 13070
rect 15182 11082 15194 13058
rect 15228 11082 15240 13058
rect 15182 11070 15240 11082
rect 15270 13058 15328 13070
rect 15270 11082 15282 13058
rect 15316 11082 15328 13058
rect 15270 11070 15328 11082
rect 15358 13058 15416 13070
rect 15358 11082 15370 13058
rect 15404 11082 15416 13058
rect 15358 11070 15416 11082
rect 15446 13058 15504 13070
rect 15446 11082 15458 13058
rect 15492 11082 15504 13058
rect 15446 11070 15504 11082
rect 15534 13058 15592 13070
rect 15534 11082 15546 13058
rect 15580 11082 15592 13058
rect 15534 11070 15592 11082
rect 15622 13058 15680 13070
rect 15622 11082 15634 13058
rect 15668 11082 15680 13058
rect 15622 11070 15680 11082
rect 15710 13058 15768 13070
rect 15710 11082 15722 13058
rect 15756 11082 15768 13058
rect 15710 11070 15768 11082
rect 15798 13058 15856 13070
rect 15798 11082 15810 13058
rect 15844 11082 15856 13058
rect 15798 11070 15856 11082
rect 15886 13058 15944 13070
rect 15886 11082 15898 13058
rect 15932 11082 15944 13058
rect 15886 11070 15944 11082
rect 15974 13058 16032 13070
rect 15974 11082 15986 13058
rect 16020 11082 16032 13058
rect 15974 11070 16032 11082
rect 16062 13058 16120 13070
rect 16062 11082 16074 13058
rect 16108 11082 16120 13058
rect 16062 11070 16120 11082
rect 16150 13058 16208 13070
rect 16150 11082 16162 13058
rect 16196 11082 16208 13058
rect 16150 11070 16208 11082
rect 16238 13058 16296 13070
rect 16238 11082 16250 13058
rect 16284 11082 16296 13058
rect 16238 11070 16296 11082
rect 16326 13058 16384 13070
rect 16326 11082 16338 13058
rect 16372 11082 16384 13058
rect 16326 11070 16384 11082
rect 16414 13058 16472 13070
rect 16414 11082 16426 13058
rect 16460 11082 16472 13058
rect 16414 11070 16472 11082
rect 16502 13058 16560 13070
rect 16502 11082 16514 13058
rect 16548 11082 16560 13058
rect 16502 11070 16560 11082
rect 16590 13058 16648 13070
rect 16590 11082 16602 13058
rect 16636 11082 16648 13058
rect 16590 11070 16648 11082
rect 16678 13058 16736 13070
rect 16678 11082 16690 13058
rect 16724 11082 16736 13058
rect 16678 11070 16736 11082
rect 16766 13058 16824 13070
rect 16766 11082 16778 13058
rect 16812 11082 16824 13058
rect 16766 11070 16824 11082
rect 16854 13058 16912 13070
rect 16854 11082 16866 13058
rect 16900 11082 16912 13058
rect 16854 11070 16912 11082
rect 16942 13058 17000 13070
rect 16942 11082 16954 13058
rect 16988 11082 17000 13058
rect 16942 11070 17000 11082
rect 17030 13058 17088 13070
rect 17030 11082 17042 13058
rect 17076 11082 17088 13058
rect 17030 11070 17088 11082
rect 17118 13058 17176 13070
rect 17118 11082 17130 13058
rect 17164 11082 17176 13058
rect 17118 11070 17176 11082
rect 17206 13058 17264 13070
rect 17206 11082 17218 13058
rect 17252 11082 17264 13058
rect 17206 11070 17264 11082
rect 17294 13058 17352 13070
rect 17294 11082 17306 13058
rect 17340 11082 17352 13058
rect 17294 11070 17352 11082
rect 17382 13058 17440 13070
rect 17382 11082 17394 13058
rect 17428 11082 17440 13058
rect 17382 11070 17440 11082
rect 17470 13058 17528 13070
rect 17470 11082 17482 13058
rect 17516 11082 17528 13058
rect 17470 11070 17528 11082
<< pdiff >>
rect 15818 23177 15880 23189
rect 15818 21201 15830 23177
rect 15864 21201 15880 23177
rect 15818 21189 15880 21201
rect 15910 23177 15976 23189
rect 15910 21201 15926 23177
rect 15960 21201 15976 23177
rect 15910 21189 15976 21201
rect 16006 23177 16072 23189
rect 16006 21201 16022 23177
rect 16056 21201 16072 23177
rect 16006 21189 16072 21201
rect 16102 23177 16164 23189
rect 16102 21201 16118 23177
rect 16152 21201 16164 23177
rect 16102 21189 16164 21201
rect 17080 15931 17142 15943
rect 17080 13955 17092 15931
rect 17126 13955 17142 15931
rect 17080 13943 17142 13955
rect 17172 15931 17238 15943
rect 17172 13955 17188 15931
rect 17222 13955 17238 15931
rect 17172 13943 17238 13955
rect 17268 15931 17334 15943
rect 17268 13955 17284 15931
rect 17318 13955 17334 15931
rect 17268 13943 17334 13955
rect 17364 15931 17426 15943
rect 17364 13955 17380 15931
rect 17414 13955 17426 15931
rect 17364 13943 17426 13955
<< ndiffc >>
rect 13970 21162 14004 23138
rect 14066 21162 14100 23138
rect 14162 21162 14196 23138
rect 14258 21162 14292 23138
rect 14354 21162 14388 23138
rect 14450 21162 14484 23138
rect 14546 21162 14580 23138
rect 14642 21162 14676 23138
rect 14738 21162 14772 23138
rect 16662 22052 16696 24028
rect 16758 22052 16792 24028
rect 16854 22052 16888 24028
rect 16950 22052 16984 24028
rect 17046 22052 17080 24028
rect 17142 22052 17176 24028
rect 17238 22052 17272 24028
rect 17334 22052 17368 24028
rect 17430 22052 17464 24028
rect 17526 22052 17560 24028
rect 17622 22052 17656 24028
rect 14830 19172 14864 20434
rect 14926 19172 14960 20434
rect 15022 19172 15056 20434
rect 15118 19172 15152 20434
rect 15214 19172 15248 20434
rect 15310 19172 15344 20434
rect 15406 19172 15440 20434
rect 15502 19172 15536 20434
rect 15990 19172 16024 19948
rect 16086 19172 16120 19948
rect 16182 19172 16216 19948
rect 16278 19172 16312 19948
rect 15016 16946 15050 18482
rect 15104 16946 15138 18482
rect 15426 16946 15460 18482
rect 15514 16946 15548 18482
rect 13572 13916 13606 15452
rect 13660 13916 13694 15452
rect 14422 13916 14456 15892
rect 14518 13916 14552 15892
rect 14614 13916 14648 15892
rect 14710 13916 14744 15892
rect 14806 13916 14840 15892
rect 14902 13916 14936 15892
rect 14998 13916 15032 15892
rect 15094 13916 15128 15892
rect 15190 13916 15224 15892
rect 13434 11082 13468 13058
rect 13522 11082 13556 13058
rect 13610 11082 13644 13058
rect 13698 11082 13732 13058
rect 13786 11082 13820 13058
rect 13874 11082 13908 13058
rect 13962 11082 13996 13058
rect 14050 11082 14084 13058
rect 14138 11082 14172 13058
rect 14226 11082 14260 13058
rect 14314 11082 14348 13058
rect 14402 11082 14436 13058
rect 14490 11082 14524 13058
rect 14578 11082 14612 13058
rect 14666 11082 14700 13058
rect 14754 11082 14788 13058
rect 14842 11082 14876 13058
rect 14930 11082 14964 13058
rect 15018 11082 15052 13058
rect 15106 11082 15140 13058
rect 15194 11082 15228 13058
rect 15282 11082 15316 13058
rect 15370 11082 15404 13058
rect 15458 11082 15492 13058
rect 15546 11082 15580 13058
rect 15634 11082 15668 13058
rect 15722 11082 15756 13058
rect 15810 11082 15844 13058
rect 15898 11082 15932 13058
rect 15986 11082 16020 13058
rect 16074 11082 16108 13058
rect 16162 11082 16196 13058
rect 16250 11082 16284 13058
rect 16338 11082 16372 13058
rect 16426 11082 16460 13058
rect 16514 11082 16548 13058
rect 16602 11082 16636 13058
rect 16690 11082 16724 13058
rect 16778 11082 16812 13058
rect 16866 11082 16900 13058
rect 16954 11082 16988 13058
rect 17042 11082 17076 13058
rect 17130 11082 17164 13058
rect 17218 11082 17252 13058
rect 17306 11082 17340 13058
rect 17394 11082 17428 13058
rect 17482 11082 17516 13058
<< pdiffc >>
rect 15830 21201 15864 23177
rect 15926 21201 15960 23177
rect 16022 21201 16056 23177
rect 16118 21201 16152 23177
rect 17092 13955 17126 15931
rect 17188 13955 17222 15931
rect 17284 13955 17318 15931
rect 17380 13955 17414 15931
<< psubdiff >>
rect 12916 24712 13012 24746
rect 16944 24712 17040 24746
rect 12916 24650 12950 24712
rect 17006 24650 17040 24712
rect 12916 24450 12950 24512
rect 17006 24450 17040 24512
rect 12916 24416 13012 24450
rect 16944 24416 17040 24450
rect 16548 24180 16644 24214
rect 17674 24180 17770 24214
rect 16548 24118 16582 24180
rect 12946 24032 13042 24066
rect 14774 24032 14870 24066
rect 12946 23970 12980 24032
rect 14836 23970 14870 24032
rect 12946 23770 12980 23832
rect 14836 23770 14870 23832
rect 12946 23736 13042 23770
rect 14774 23736 14870 23770
rect 15176 23326 15272 23360
rect 15410 23326 15506 23360
rect 13856 23290 13952 23324
rect 14790 23290 14886 23324
rect 13856 23228 13890 23290
rect 13356 22166 13452 22200
rect 13590 22166 13686 22200
rect 13356 22104 13390 22166
rect 13652 22104 13686 22166
rect 13356 21010 13390 21072
rect 13652 21010 13686 21072
rect 13356 20976 13452 21010
rect 13590 20976 13686 21010
rect 14852 23228 14886 23290
rect 13856 21010 13890 21072
rect 14852 21010 14886 21072
rect 13856 20976 13952 21010
rect 14790 20976 14886 21010
rect 15176 23264 15210 23326
rect 15472 23264 15506 23326
rect 15176 21030 15210 21092
rect 15472 21030 15506 21092
rect 15176 20996 15272 21030
rect 15410 20996 15506 21030
rect 17736 24118 17770 24180
rect 16548 21900 16582 21962
rect 17736 21900 17770 21962
rect 16548 21866 16644 21900
rect 17674 21866 17770 21900
rect 16656 21446 16752 21480
rect 16890 21446 16986 21480
rect 16656 21384 16690 21446
rect 14716 20586 14812 20620
rect 15554 20586 15650 20620
rect 14716 20524 14750 20586
rect 13182 19826 13278 19860
rect 14348 19826 14444 19860
rect 13182 19764 13216 19826
rect 14410 19764 14444 19826
rect 13182 16794 13216 16856
rect 15616 20524 15650 20586
rect 14716 19020 14750 19082
rect 15616 19020 15650 19082
rect 14716 18986 14812 19020
rect 15554 18986 15650 19020
rect 15876 20100 15972 20134
rect 16330 20100 16426 20134
rect 15876 20038 15910 20100
rect 16392 20038 16426 20100
rect 15876 19020 15910 19082
rect 16392 19020 16426 19082
rect 15876 18986 15972 19020
rect 16330 18986 16426 19020
rect 16952 21384 16986 21446
rect 16656 18790 16690 18852
rect 16952 18790 16986 18852
rect 16656 18756 16752 18790
rect 16890 18756 16986 18790
rect 17266 21466 17362 21500
rect 17500 21466 17596 21500
rect 17266 21404 17300 21466
rect 14902 18634 14998 18668
rect 15156 18634 15252 18668
rect 14902 18572 14936 18634
rect 14410 16794 14444 16856
rect 13182 16760 13278 16794
rect 14348 16760 14444 16794
rect 14512 17950 14608 17984
rect 14746 17950 14842 17984
rect 14512 17888 14546 17950
rect 14808 17888 14842 17950
rect 14512 16794 14546 16856
rect 14808 16794 14842 16856
rect 14512 16760 14608 16794
rect 14746 16760 14842 16794
rect 15218 18572 15252 18634
rect 14902 16794 14936 16856
rect 15218 16794 15252 16856
rect 14902 16760 14998 16794
rect 15156 16760 15252 16794
rect 15312 18634 15408 18668
rect 15566 18634 15662 18668
rect 15312 18572 15346 18634
rect 15628 18572 15662 18634
rect 15312 16794 15346 16856
rect 16124 18651 16220 18685
rect 16358 18651 16454 18685
rect 16124 18589 16158 18651
rect 15628 16794 15662 16856
rect 15312 16760 15408 16794
rect 15566 16760 15662 16794
rect 15732 17950 15828 17984
rect 15966 17950 16062 17984
rect 15732 17888 15766 17950
rect 16028 17888 16062 17950
rect 15732 16794 15766 16856
rect 16028 16794 16062 16856
rect 15732 16760 15828 16794
rect 15966 16760 16062 16794
rect 16420 18589 16454 18651
rect 16124 16795 16158 16857
rect 16686 18426 16782 18460
rect 16884 18426 16980 18460
rect 16686 18364 16720 18426
rect 16946 18364 16980 18426
rect 16686 18200 16720 18262
rect 16946 18200 16980 18262
rect 16686 18166 16782 18200
rect 16884 18166 16980 18200
rect 17562 21404 17596 21466
rect 17266 17410 17300 17472
rect 17562 17410 17596 17472
rect 17266 17376 17362 17410
rect 17500 17376 17596 17410
rect 16420 16795 16454 16857
rect 16124 16761 16220 16795
rect 16358 16761 16454 16795
rect 14308 16044 14404 16078
rect 15242 16044 15338 16078
rect 14308 15982 14342 16044
rect 13458 15604 13554 15638
rect 13712 15604 13808 15638
rect 13458 15542 13492 15604
rect 13774 15542 13808 15604
rect 13458 13764 13492 13826
rect 13774 13764 13808 13826
rect 13458 13730 13554 13764
rect 13712 13730 13808 13764
rect 15304 15982 15338 16044
rect 14308 13764 14342 13826
rect 15304 13764 15338 13826
rect 14308 13730 14404 13764
rect 15242 13730 15338 13764
rect 16018 16060 16114 16094
rect 16252 16060 16348 16094
rect 16018 15998 16052 16060
rect 16314 15998 16348 16060
rect 16018 13764 16052 13826
rect 16314 13764 16348 13826
rect 16018 13730 16114 13764
rect 16252 13730 16348 13764
rect 13074 13571 17870 13590
rect 13074 13488 13313 13571
rect 17596 13488 17870 13571
rect 13074 13455 17870 13488
rect 13074 13424 13209 13455
rect 13074 10790 13103 13424
rect 13176 10790 13209 13424
rect 17728 13433 17870 13455
rect 13074 10738 13209 10790
rect 17728 10799 17766 13433
rect 17839 10799 17870 13433
rect 17728 10738 17870 10799
rect 13074 10718 17870 10738
rect 13074 10635 13355 10718
rect 17638 10635 17870 10718
rect 13074 10610 17870 10635
<< nsubdiff >>
rect 15716 23338 15812 23372
rect 16170 23338 16266 23372
rect 15716 23276 15750 23338
rect 16232 23276 16266 23338
rect 15716 21040 15750 21102
rect 16232 21040 16266 21102
rect 15716 21006 15812 21040
rect 16170 21006 16266 21040
rect 16978 16092 17074 16126
rect 17432 16092 17528 16126
rect 16978 16030 17012 16092
rect 17494 16030 17528 16092
rect 16978 13794 17012 13856
rect 17494 13794 17528 13856
rect 16978 13760 17074 13794
rect 17432 13760 17528 13794
<< psubdiffcont >>
rect 13012 24712 16944 24746
rect 12916 24512 12950 24650
rect 17006 24512 17040 24650
rect 13012 24416 16944 24450
rect 16644 24180 17674 24214
rect 13042 24032 14774 24066
rect 12946 23832 12980 23970
rect 14836 23832 14870 23970
rect 13042 23736 14774 23770
rect 15272 23326 15410 23360
rect 13952 23290 14790 23324
rect 13452 22166 13590 22200
rect 13356 21072 13390 22104
rect 13652 21072 13686 22104
rect 13452 20976 13590 21010
rect 13856 21072 13890 23228
rect 14852 21072 14886 23228
rect 13952 20976 14790 21010
rect 15176 21092 15210 23264
rect 15472 21092 15506 23264
rect 15272 20996 15410 21030
rect 16548 21962 16582 24118
rect 17736 21962 17770 24118
rect 16644 21866 17674 21900
rect 16752 21446 16890 21480
rect 14812 20586 15554 20620
rect 13278 19826 14348 19860
rect 13182 16856 13216 19764
rect 14410 16856 14444 19764
rect 14716 19082 14750 20524
rect 15616 19082 15650 20524
rect 14812 18986 15554 19020
rect 15972 20100 16330 20134
rect 15876 19082 15910 20038
rect 16392 19082 16426 20038
rect 15972 18986 16330 19020
rect 16656 18852 16690 21384
rect 16952 18852 16986 21384
rect 16752 18756 16890 18790
rect 17362 21466 17500 21500
rect 14998 18634 15156 18668
rect 13278 16760 14348 16794
rect 14608 17950 14746 17984
rect 14512 16856 14546 17888
rect 14808 16856 14842 17888
rect 14608 16760 14746 16794
rect 14902 16856 14936 18572
rect 15218 16856 15252 18572
rect 14998 16760 15156 16794
rect 15408 18634 15566 18668
rect 15312 16856 15346 18572
rect 15628 16856 15662 18572
rect 16220 18651 16358 18685
rect 15408 16760 15566 16794
rect 15828 17950 15966 17984
rect 15732 16856 15766 17888
rect 16028 16856 16062 17888
rect 15828 16760 15966 16794
rect 16124 16857 16158 18589
rect 16420 16857 16454 18589
rect 16782 18426 16884 18460
rect 16686 18262 16720 18364
rect 16946 18262 16980 18364
rect 16782 18166 16884 18200
rect 17266 17472 17300 21404
rect 17562 17472 17596 21404
rect 17362 17376 17500 17410
rect 16220 16761 16358 16795
rect 14404 16044 15242 16078
rect 13554 15604 13712 15638
rect 13458 13826 13492 15542
rect 13774 13826 13808 15542
rect 13554 13730 13712 13764
rect 14308 13826 14342 15982
rect 15304 13826 15338 15982
rect 14404 13730 15242 13764
rect 16114 16060 16252 16094
rect 16018 13826 16052 15998
rect 16314 13826 16348 15998
rect 16114 13730 16252 13764
rect 13313 13488 17596 13571
rect 13103 10790 13176 13424
rect 17766 10799 17839 13433
rect 13355 10635 17638 10718
<< nsubdiffcont >>
rect 15812 23338 16170 23372
rect 15716 21102 15750 23276
rect 16232 21102 16266 23276
rect 15812 21006 16170 21040
rect 17074 16092 17432 16126
rect 16978 13856 17012 16030
rect 17494 13856 17528 16030
rect 17074 13760 17432 13794
<< poly >>
rect 14020 23222 14164 23238
rect 14020 23188 14114 23222
rect 14148 23188 14164 23222
rect 14020 23172 14164 23188
rect 14290 23222 14356 23238
rect 14290 23188 14306 23222
rect 14340 23188 14356 23222
rect 14020 23150 14050 23172
rect 14116 23150 14146 23172
rect 14212 23150 14242 23176
rect 14290 23172 14356 23188
rect 14482 23222 14548 23238
rect 14482 23188 14498 23222
rect 14532 23188 14548 23222
rect 14308 23150 14338 23172
rect 14404 23150 14434 23176
rect 14482 23172 14548 23188
rect 14674 23222 14740 23238
rect 14674 23188 14690 23222
rect 14724 23188 14740 23222
rect 14500 23150 14530 23172
rect 14596 23150 14626 23176
rect 14674 23172 14740 23188
rect 14692 23150 14722 23172
rect 14020 21128 14050 21150
rect 14002 21112 14068 21128
rect 14116 21124 14146 21150
rect 14212 21128 14242 21150
rect 14002 21078 14018 21112
rect 14052 21078 14068 21112
rect 14002 21062 14068 21078
rect 14194 21112 14260 21128
rect 14308 21124 14338 21150
rect 14404 21128 14434 21150
rect 14194 21078 14210 21112
rect 14244 21078 14260 21112
rect 14194 21062 14260 21078
rect 14386 21112 14452 21128
rect 14500 21124 14530 21150
rect 14596 21128 14626 21150
rect 14692 21128 14722 21150
rect 14386 21078 14402 21112
rect 14436 21078 14452 21112
rect 14386 21062 14452 21078
rect 14578 21112 14722 21128
rect 14578 21078 14594 21112
rect 14628 21078 14722 21112
rect 14578 21062 14722 21078
rect 15958 23270 16024 23286
rect 15958 23236 15974 23270
rect 16008 23236 16024 23270
rect 15958 23220 16024 23236
rect 15880 23189 15910 23215
rect 15976 23189 16006 23220
rect 16072 23189 16102 23215
rect 15880 21160 15910 21189
rect 15976 21160 16006 21189
rect 16072 21160 16102 21189
rect 15861 21142 16120 21160
rect 15861 21108 15878 21142
rect 15912 21108 16070 21142
rect 16104 21108 16120 21142
rect 15861 21091 16120 21108
rect 16710 24112 16860 24130
rect 16710 24078 16806 24112
rect 16840 24078 16860 24112
rect 16710 24060 16860 24078
rect 16982 24112 17048 24128
rect 16982 24078 16998 24112
rect 17032 24078 17048 24112
rect 16712 24040 16742 24060
rect 16808 24040 16838 24060
rect 16904 24040 16934 24066
rect 16982 24062 17048 24078
rect 17174 24112 17240 24128
rect 17174 24078 17190 24112
rect 17224 24078 17240 24112
rect 17000 24040 17030 24062
rect 17096 24040 17126 24066
rect 17174 24062 17240 24078
rect 17366 24112 17432 24128
rect 17366 24078 17382 24112
rect 17416 24078 17432 24112
rect 17192 24040 17222 24062
rect 17288 24040 17318 24066
rect 17366 24062 17432 24078
rect 17558 24112 17624 24128
rect 17558 24078 17574 24112
rect 17608 24078 17624 24112
rect 17384 24040 17414 24062
rect 17480 24040 17510 24066
rect 17558 24062 17624 24078
rect 17576 24040 17606 24062
rect 16712 22018 16742 22040
rect 16694 22002 16760 22018
rect 16808 22014 16838 22040
rect 16904 22018 16934 22040
rect 16694 21968 16710 22002
rect 16744 21968 16760 22002
rect 16694 21952 16760 21968
rect 16886 22002 16952 22018
rect 17000 22014 17030 22040
rect 17096 22018 17126 22040
rect 16886 21968 16902 22002
rect 16936 21968 16952 22002
rect 16886 21952 16952 21968
rect 17078 22002 17144 22018
rect 17192 22014 17222 22040
rect 17288 22018 17318 22040
rect 17078 21968 17094 22002
rect 17128 21968 17144 22002
rect 17078 21952 17144 21968
rect 17270 22002 17336 22018
rect 17384 22014 17414 22040
rect 17480 22020 17510 22040
rect 17576 22020 17606 22040
rect 17270 21968 17286 22002
rect 17320 21968 17336 22002
rect 17270 21952 17336 21968
rect 17460 22002 17610 22020
rect 17460 21968 17478 22002
rect 17512 21968 17610 22002
rect 17460 21950 17610 21968
rect 14880 20518 15490 20540
rect 14880 20484 14974 20518
rect 15008 20484 15166 20518
rect 15200 20484 15358 20518
rect 15392 20484 15490 20518
rect 14880 20470 15490 20484
rect 14880 20446 14910 20470
rect 14958 20468 15024 20470
rect 14976 20446 15006 20468
rect 15072 20446 15102 20470
rect 15150 20468 15216 20470
rect 15168 20446 15198 20468
rect 15264 20446 15294 20470
rect 15342 20468 15408 20470
rect 15360 20446 15390 20468
rect 15456 20446 15486 20470
rect 14880 19140 14910 19160
rect 14976 19140 15006 19160
rect 15072 19140 15102 19160
rect 15168 19140 15198 19160
rect 15264 19140 15294 19160
rect 15360 19140 15390 19160
rect 15456 19140 15486 19160
rect 14860 19122 15510 19140
rect 14860 19088 14878 19122
rect 14912 19088 15070 19122
rect 15104 19088 15262 19122
rect 15296 19088 15454 19122
rect 15488 19088 15510 19122
rect 14860 19070 15510 19088
rect 16040 20032 16270 20050
rect 16040 19998 16134 20032
rect 16168 19998 16270 20032
rect 16040 19980 16270 19998
rect 16040 19960 16070 19980
rect 16136 19960 16166 19980
rect 16232 19960 16262 19980
rect 16040 19140 16070 19160
rect 16136 19140 16166 19160
rect 16232 19140 16262 19160
rect 16020 19122 16280 19140
rect 16020 19088 16038 19122
rect 16072 19088 16230 19122
rect 16264 19088 16280 19122
rect 16020 19070 16280 19088
rect 15044 18566 15110 18582
rect 15044 18532 15060 18566
rect 15094 18532 15110 18566
rect 15044 18516 15110 18532
rect 15062 18494 15092 18516
rect 15062 16912 15092 16934
rect 15044 16896 15110 16912
rect 15044 16862 15060 16896
rect 15094 16862 15110 16896
rect 15044 16846 15110 16862
rect 15454 18566 15520 18582
rect 15454 18532 15470 18566
rect 15504 18532 15520 18566
rect 15454 18516 15520 18532
rect 15472 18494 15502 18516
rect 15472 16912 15502 16934
rect 15454 16896 15520 16912
rect 15454 16862 15470 16896
rect 15504 16862 15520 16896
rect 15454 16846 15520 16862
rect 13598 15536 13666 15554
rect 13598 15502 13616 15536
rect 13650 15502 13666 15536
rect 13598 15496 13666 15502
rect 13600 15486 13666 15496
rect 13618 15464 13648 15486
rect 13618 13882 13648 13904
rect 13600 13866 13666 13882
rect 13600 13832 13616 13866
rect 13650 13832 13666 13866
rect 13600 13816 13666 13832
rect 14472 15976 14622 15994
rect 14472 15942 14566 15976
rect 14600 15942 14622 15976
rect 14472 15924 14622 15942
rect 14742 15976 14808 15992
rect 14742 15942 14758 15976
rect 14792 15942 14808 15976
rect 14472 15904 14502 15924
rect 14568 15904 14598 15924
rect 14664 15904 14694 15930
rect 14742 15926 14808 15942
rect 14934 15976 15000 15992
rect 14934 15942 14950 15976
rect 14984 15942 15000 15976
rect 14760 15904 14790 15926
rect 14856 15904 14886 15930
rect 14934 15926 15000 15942
rect 15126 15976 15192 15992
rect 15126 15942 15142 15976
rect 15176 15942 15192 15976
rect 14952 15904 14982 15926
rect 15048 15904 15078 15930
rect 15126 15926 15192 15942
rect 15144 15904 15174 15926
rect 14472 13882 14502 13904
rect 14454 13866 14520 13882
rect 14568 13878 14598 13904
rect 14664 13882 14694 13904
rect 14454 13832 14470 13866
rect 14504 13832 14520 13866
rect 14454 13816 14520 13832
rect 14646 13866 14712 13882
rect 14760 13878 14790 13904
rect 14856 13882 14886 13904
rect 14646 13832 14662 13866
rect 14696 13832 14712 13866
rect 14646 13816 14712 13832
rect 14838 13866 14904 13882
rect 14952 13878 14982 13904
rect 15048 13882 15078 13904
rect 15144 13882 15174 13904
rect 14838 13832 14854 13866
rect 14888 13832 14904 13866
rect 14838 13816 14904 13832
rect 15030 13866 15174 13882
rect 15030 13832 15046 13866
rect 15080 13832 15174 13866
rect 15030 13816 15174 13832
rect 17142 16024 17364 16040
rect 17142 15990 17236 16024
rect 17270 15990 17364 16024
rect 17142 15969 17364 15990
rect 17142 15943 17172 15969
rect 17238 15943 17268 15969
rect 17334 15943 17364 15969
rect 17142 13917 17172 13943
rect 17238 13917 17268 13943
rect 17334 13917 17364 13943
rect 17124 13896 17382 13917
rect 17124 13862 17140 13896
rect 17174 13862 17332 13896
rect 17366 13862 17382 13896
rect 17124 13846 17382 13862
rect 17000 13313 17118 13334
rect 17000 13273 17021 13313
rect 17093 13273 17118 13313
rect 17000 13254 17118 13273
rect 13480 13195 13571 13215
rect 13480 13133 13500 13195
rect 13552 13175 13571 13195
rect 13675 13177 13750 13195
rect 13552 13133 13598 13175
rect 13675 13172 13689 13177
rect 13480 13096 13598 13133
rect 13480 13070 13510 13096
rect 13568 13070 13598 13096
rect 13656 13131 13689 13172
rect 13736 13172 13750 13177
rect 14029 13173 14104 13191
rect 13736 13131 13774 13172
rect 14029 13170 14043 13173
rect 13656 13115 13774 13131
rect 13656 13070 13686 13115
rect 13744 13070 13774 13115
rect 14008 13127 14043 13170
rect 14090 13170 14104 13173
rect 14382 13172 14457 13189
rect 14735 13172 14810 13190
rect 15086 13172 15161 13190
rect 15440 13173 15515 13191
rect 15790 13173 15865 13190
rect 15440 13172 15454 13173
rect 14360 13171 14478 13172
rect 14090 13127 14126 13170
rect 14008 13111 14126 13127
rect 13832 13070 13862 13096
rect 13920 13070 13950 13096
rect 14008 13070 14038 13111
rect 14096 13070 14126 13111
rect 14360 13125 14396 13171
rect 14443 13125 14478 13171
rect 14360 13109 14478 13125
rect 14184 13070 14214 13096
rect 14272 13070 14302 13096
rect 14360 13070 14390 13109
rect 14448 13070 14478 13109
rect 14712 13126 14749 13172
rect 14796 13126 14830 13172
rect 14712 13110 14830 13126
rect 14536 13070 14566 13096
rect 14624 13070 14654 13096
rect 14712 13070 14742 13110
rect 14800 13070 14830 13110
rect 15064 13126 15100 13172
rect 15147 13126 15182 13172
rect 15064 13110 15182 13126
rect 14888 13070 14918 13096
rect 14976 13070 15006 13096
rect 15064 13070 15094 13110
rect 15152 13070 15182 13110
rect 15416 13127 15454 13172
rect 15501 13172 15515 13173
rect 15768 13172 15886 13173
rect 16142 13172 16217 13189
rect 16495 13172 16570 13189
rect 16844 13172 16919 13189
rect 15501 13127 15534 13172
rect 15416 13111 15534 13127
rect 15240 13070 15270 13096
rect 15328 13070 15358 13096
rect 15416 13070 15446 13111
rect 15504 13070 15534 13111
rect 15768 13126 15804 13172
rect 15851 13126 15886 13172
rect 15768 13110 15886 13126
rect 15592 13070 15622 13096
rect 15680 13070 15710 13096
rect 15768 13070 15798 13110
rect 15856 13070 15886 13110
rect 16120 13171 16238 13172
rect 16120 13125 16156 13171
rect 16203 13125 16238 13171
rect 16120 13109 16238 13125
rect 15944 13070 15974 13096
rect 16032 13070 16062 13096
rect 16120 13070 16150 13109
rect 16208 13070 16238 13109
rect 16472 13171 16590 13172
rect 16472 13125 16509 13171
rect 16556 13125 16590 13171
rect 16472 13109 16590 13125
rect 16296 13070 16326 13096
rect 16384 13070 16414 13096
rect 16472 13070 16502 13109
rect 16560 13070 16590 13109
rect 16824 13171 16942 13172
rect 16824 13125 16858 13171
rect 16905 13125 16942 13171
rect 16824 13109 16942 13125
rect 16648 13070 16678 13096
rect 16736 13070 16766 13096
rect 16824 13070 16854 13109
rect 16912 13070 16942 13109
rect 17000 13070 17030 13254
rect 17088 13070 17118 13254
rect 17198 13173 17273 13189
rect 17176 13171 17294 13173
rect 17176 13125 17212 13171
rect 17259 13125 17294 13171
rect 17371 13171 17446 13189
rect 17371 13164 17385 13171
rect 17176 13109 17294 13125
rect 17176 13070 17206 13109
rect 17264 13070 17294 13109
rect 17352 13125 17385 13164
rect 17432 13164 17446 13171
rect 17432 13125 17470 13164
rect 17352 13109 17470 13125
rect 17352 13070 17382 13109
rect 17440 13070 17470 13109
rect 13480 11020 13510 11070
rect 13568 11020 13598 11070
rect 13656 11044 13686 11070
rect 13744 11044 13774 11070
rect 13480 11002 13598 11020
rect 13480 10970 13511 11002
rect 13497 10956 13511 10970
rect 13558 10970 13598 11002
rect 13832 11014 13862 11070
rect 13920 11014 13950 11070
rect 14008 11044 14038 11070
rect 14096 11044 14126 11070
rect 13832 10996 13950 11014
rect 13558 10956 13572 10970
rect 13832 10969 13861 10996
rect 13497 10940 13572 10956
rect 13847 10950 13861 10969
rect 13908 10969 13950 10996
rect 14184 11017 14214 11070
rect 14272 11017 14302 11070
rect 14360 11044 14390 11070
rect 14448 11044 14478 11070
rect 14184 10999 14302 11017
rect 14184 10969 14219 10999
rect 13908 10950 13922 10969
rect 13847 10934 13922 10950
rect 14205 10953 14219 10969
rect 14266 10969 14302 10999
rect 14536 11017 14566 11070
rect 14624 11017 14654 11070
rect 14712 11044 14742 11070
rect 14800 11044 14830 11070
rect 14536 10999 14654 11017
rect 14536 10969 14567 10999
rect 14266 10953 14280 10969
rect 14205 10937 14280 10953
rect 14553 10953 14567 10969
rect 14614 10969 14654 10999
rect 14888 11017 14918 11070
rect 14976 11017 15006 11070
rect 15064 11044 15094 11070
rect 15152 11044 15182 11070
rect 14888 10999 15006 11017
rect 14888 10970 14918 10999
rect 14614 10953 14628 10969
rect 14553 10937 14628 10953
rect 14904 10953 14918 10970
rect 14965 10970 15006 10999
rect 15240 11016 15270 11070
rect 15328 11016 15358 11070
rect 15416 11044 15446 11070
rect 15504 11044 15534 11070
rect 15240 10998 15358 11016
rect 15240 10970 15269 10998
rect 14965 10953 14979 10970
rect 14904 10937 14979 10953
rect 15255 10952 15269 10970
rect 15316 10970 15358 10998
rect 15592 11014 15622 11070
rect 15680 11014 15710 11070
rect 15768 11044 15798 11070
rect 15856 11044 15886 11070
rect 15592 10996 15710 11014
rect 15592 10971 15620 10996
rect 15316 10952 15330 10970
rect 15255 10936 15330 10952
rect 15606 10950 15620 10971
rect 15667 10971 15710 10996
rect 15944 11017 15974 11070
rect 16032 11017 16062 11070
rect 16120 11044 16150 11070
rect 16208 11044 16238 11070
rect 15944 10999 16062 11017
rect 15944 10971 15975 10999
rect 15667 10950 15681 10971
rect 15606 10934 15681 10950
rect 15961 10953 15975 10971
rect 16022 10971 16062 10999
rect 16296 11013 16326 11070
rect 16384 11013 16414 11070
rect 16472 11044 16502 11070
rect 16560 11044 16590 11070
rect 16296 10995 16414 11013
rect 16296 10971 16325 10995
rect 16022 10953 16036 10971
rect 15961 10937 16036 10953
rect 16311 10949 16325 10971
rect 16372 10971 16414 10995
rect 16648 11015 16678 11070
rect 16736 11015 16766 11070
rect 16824 11044 16854 11070
rect 16912 11044 16942 11070
rect 16648 10997 16766 11015
rect 16372 10949 16386 10971
rect 16648 10970 16679 10997
rect 16311 10933 16386 10949
rect 16665 10951 16679 10970
rect 16726 10970 16766 10997
rect 17000 11013 17030 11070
rect 17088 11013 17118 11070
rect 17176 11044 17206 11070
rect 17264 11044 17294 11070
rect 17000 10995 17118 11013
rect 17000 10971 17029 10995
rect 16726 10951 16740 10970
rect 16665 10935 16740 10951
rect 17015 10949 17029 10971
rect 17076 10971 17118 10995
rect 17352 11024 17382 11070
rect 17440 11024 17470 11070
rect 17352 10994 17472 11024
rect 17076 10949 17090 10971
rect 17015 10933 17090 10949
rect 17352 10914 17372 10994
rect 17452 10914 17472 10994
rect 17352 10884 17472 10914
<< polycont >>
rect 14114 23188 14148 23222
rect 14306 23188 14340 23222
rect 14498 23188 14532 23222
rect 14690 23188 14724 23222
rect 14018 21078 14052 21112
rect 14210 21078 14244 21112
rect 14402 21078 14436 21112
rect 14594 21078 14628 21112
rect 15974 23236 16008 23270
rect 15878 21108 15912 21142
rect 16070 21108 16104 21142
rect 16806 24078 16840 24112
rect 16998 24078 17032 24112
rect 17190 24078 17224 24112
rect 17382 24078 17416 24112
rect 17574 24078 17608 24112
rect 16710 21968 16744 22002
rect 16902 21968 16936 22002
rect 17094 21968 17128 22002
rect 17286 21968 17320 22002
rect 17478 21968 17512 22002
rect 14974 20484 15008 20518
rect 15166 20484 15200 20518
rect 15358 20484 15392 20518
rect 14878 19088 14912 19122
rect 15070 19088 15104 19122
rect 15262 19088 15296 19122
rect 15454 19088 15488 19122
rect 16134 19998 16168 20032
rect 16038 19088 16072 19122
rect 16230 19088 16264 19122
rect 15060 18532 15094 18566
rect 15060 16862 15094 16896
rect 15470 18532 15504 18566
rect 15470 16862 15504 16896
rect 13616 15502 13650 15536
rect 13616 13832 13650 13866
rect 14566 15942 14600 15976
rect 14758 15942 14792 15976
rect 14950 15942 14984 15976
rect 15142 15942 15176 15976
rect 14470 13832 14504 13866
rect 14662 13832 14696 13866
rect 14854 13832 14888 13866
rect 15046 13832 15080 13866
rect 17236 15990 17270 16024
rect 17140 13862 17174 13896
rect 17332 13862 17366 13896
rect 17021 13273 17093 13313
rect 13500 13133 13552 13195
rect 13689 13131 13736 13177
rect 14043 13127 14090 13173
rect 14396 13125 14443 13171
rect 14749 13126 14796 13172
rect 15100 13126 15147 13172
rect 15454 13127 15501 13173
rect 15804 13126 15851 13172
rect 16156 13125 16203 13171
rect 16509 13125 16556 13171
rect 16858 13125 16905 13171
rect 17212 13125 17259 13171
rect 17385 13125 17432 13171
rect 13511 10956 13558 11002
rect 13861 10950 13908 10996
rect 14219 10953 14266 10999
rect 14567 10953 14614 10999
rect 14918 10953 14965 10999
rect 15269 10952 15316 10998
rect 15620 10950 15667 10996
rect 15975 10953 16022 10999
rect 16325 10949 16372 10995
rect 16679 10951 16726 10997
rect 17029 10949 17076 10995
rect 17372 10914 17452 10994
<< xpolycontact >>
rect 13046 24546 13478 24616
rect 16478 24546 16910 24616
rect 13076 23866 13508 23936
rect 14308 23866 14740 23936
rect 13486 21638 13556 22070
rect 13486 21106 13556 21538
rect 15306 22798 15376 23230
rect 15306 21126 15376 21558
rect 13312 19592 13744 19730
rect 13882 19592 14314 19730
rect 13312 19206 13744 19344
rect 13882 19206 14314 19344
rect 13312 18820 13744 18958
rect 13882 18820 14314 18958
rect 13312 18434 13744 18572
rect 13882 18434 14314 18572
rect 13312 18048 13744 18186
rect 13882 18048 14314 18186
rect 13312 17662 13744 17800
rect 13882 17662 14314 17800
rect 13312 17276 13744 17414
rect 13882 17276 14314 17414
rect 13312 16890 13744 17028
rect 13882 16890 14314 17028
rect 16786 20918 16856 21350
rect 16786 18886 16856 19318
rect 14642 17422 14712 17854
rect 14642 16890 14712 17322
rect 15862 17422 15932 17854
rect 15862 16890 15932 17322
rect 16254 18123 16324 18555
rect 16254 16891 16324 17323
rect 17396 20938 17466 21370
rect 17396 17506 17466 17938
rect 16148 15532 16218 15964
rect 16148 13860 16218 14292
<< ppolyres >>
rect 13478 24546 16478 24616
rect 13508 23866 14308 23936
rect 13486 21538 13556 21638
rect 15306 21558 15376 22798
rect 13744 19592 13882 19730
rect 13744 19206 13882 19344
rect 13744 18820 13882 18958
rect 13744 18434 13882 18572
rect 13744 18048 13882 18186
rect 13744 17662 13882 17800
rect 13744 17276 13882 17414
rect 13744 16890 13882 17028
rect 16786 19318 16856 20918
rect 14642 17322 14712 17422
rect 15862 17322 15932 17422
rect 16254 17323 16324 18123
rect 17396 17938 17466 20938
rect 16148 14292 16218 15532
<< ndiode >>
rect 16788 18346 16878 18358
rect 16788 18280 16800 18346
rect 16866 18280 16878 18346
rect 16788 18268 16878 18280
<< ndiodec >>
rect 16800 18280 16866 18346
<< locali >>
rect 14004 28832 16526 28932
rect 14004 27684 14118 28832
rect 16404 27684 16526 28832
rect 14004 25334 16526 27684
rect 12670 24852 17790 25334
rect 12670 23542 12834 24852
rect 13049 24746 13484 24749
rect 12916 24712 13012 24746
rect 16944 24712 17040 24746
rect 12916 24650 12950 24712
rect 13049 24616 13484 24712
rect 17006 24650 17040 24712
rect 13478 24546 13484 24616
rect 13049 24541 13484 24546
rect 12916 24450 12950 24512
rect 17006 24450 17040 24512
rect 12916 24416 13012 24450
rect 16944 24416 17040 24450
rect 16548 24180 16644 24214
rect 17674 24180 17770 24214
rect 16548 24118 16582 24180
rect 12946 24032 13042 24066
rect 14774 24032 14870 24066
rect 12946 23970 12980 24032
rect 14836 23970 14870 24032
rect 12946 23770 12980 23832
rect 14836 23770 14870 23832
rect 12946 23736 13042 23770
rect 14774 23736 14870 23770
rect 13300 23580 15938 23584
rect 12926 23579 15938 23580
rect 16270 23579 16450 23580
rect 12926 23560 16450 23579
rect 12926 23550 16290 23560
rect 12926 23542 13090 23550
rect 12670 23390 13090 23542
rect 13310 23430 16290 23550
rect 16430 23430 16450 23560
rect 13310 23414 16450 23430
rect 12670 23378 13310 23390
rect 12926 23372 13310 23378
rect 15709 23410 16450 23414
rect 15709 23372 16448 23410
rect 15176 23326 15272 23360
rect 15410 23326 15506 23360
rect 15709 23338 15812 23372
rect 16170 23338 16448 23372
rect 15709 23332 16448 23338
rect 13856 23290 13952 23324
rect 14790 23290 14886 23324
rect 13856 23228 13890 23290
rect 13356 22166 13452 22200
rect 13590 22166 13686 22200
rect 13356 22104 13390 22166
rect 13652 22104 13686 22166
rect 13356 21010 13390 21072
rect 13652 21010 13686 21072
rect 13356 20976 13452 21010
rect 13590 20976 13686 21010
rect 14852 23228 14886 23290
rect 14098 23188 14114 23222
rect 14148 23188 14164 23222
rect 14290 23188 14306 23222
rect 14340 23188 14356 23222
rect 14482 23188 14498 23222
rect 14532 23188 14548 23222
rect 14674 23188 14690 23222
rect 14724 23188 14740 23222
rect 13970 23138 14004 23154
rect 13970 21146 14004 21162
rect 14066 23138 14100 23154
rect 14066 21146 14100 21162
rect 14162 23138 14196 23154
rect 14162 21146 14196 21162
rect 14258 23138 14292 23154
rect 14258 21146 14292 21162
rect 14354 23138 14388 23154
rect 14354 21146 14388 21162
rect 14450 23138 14484 23154
rect 14450 21146 14484 21162
rect 14546 23138 14580 23154
rect 14546 21146 14580 21162
rect 14642 23138 14676 23154
rect 14642 21146 14676 21162
rect 14738 23138 14772 23154
rect 14820 23140 14852 23150
rect 15176 23264 15210 23326
rect 14886 23140 14910 23150
rect 14820 23040 14830 23140
rect 14900 23040 14910 23140
rect 14820 23030 14852 23040
rect 14738 21146 14772 21162
rect 14002 21078 14018 21112
rect 14052 21078 14068 21112
rect 14194 21078 14210 21112
rect 14244 21078 14260 21112
rect 14386 21078 14402 21112
rect 14436 21078 14452 21112
rect 14578 21078 14594 21112
rect 14628 21078 14644 21112
rect 13856 21010 13890 21072
rect 14886 23030 14910 23040
rect 14852 21010 14886 21072
rect 13856 20976 13952 21010
rect 14790 20976 14886 21010
rect 15472 23264 15506 23326
rect 15176 21030 15210 21092
rect 15472 21030 15506 21092
rect 15176 20996 15272 21030
rect 15410 20996 15506 21030
rect 15716 23276 15750 23332
rect 16232 23276 16266 23332
rect 15958 23236 15974 23270
rect 16008 23236 16024 23270
rect 15830 23177 15864 23193
rect 15830 21185 15864 21201
rect 15926 23177 15960 23193
rect 15926 21185 15960 21201
rect 16022 23177 16056 23193
rect 16022 21185 16056 21201
rect 16118 23190 16152 23193
rect 16118 23177 16232 23190
rect 16152 23070 16232 23177
rect 16225 21565 16232 21775
rect 16118 21185 16152 21201
rect 15862 21108 15878 21142
rect 15912 21108 15928 21142
rect 16054 21108 16070 21142
rect 16104 21108 16120 21142
rect 15716 21040 15750 21102
rect 16266 23070 16270 23190
rect 17736 24118 17770 24180
rect 16790 24078 16806 24112
rect 16840 24078 16856 24112
rect 16982 24078 16998 24112
rect 17032 24078 17048 24112
rect 17174 24078 17190 24112
rect 17224 24078 17240 24112
rect 17366 24078 17382 24112
rect 17416 24078 17432 24112
rect 17558 24078 17574 24112
rect 17608 24078 17624 24112
rect 16662 24028 16696 24044
rect 16662 22036 16696 22052
rect 16758 24028 16792 24044
rect 16758 22036 16792 22052
rect 16854 24028 16888 24044
rect 16854 22036 16888 22052
rect 16950 24028 16984 24044
rect 16950 22036 16984 22052
rect 17046 24028 17080 24044
rect 17046 22036 17080 22052
rect 17142 24028 17176 24044
rect 17142 22036 17176 22052
rect 17238 24028 17272 24044
rect 17238 22036 17272 22052
rect 17334 24028 17368 24044
rect 17334 22036 17368 22052
rect 17430 24028 17464 24044
rect 17430 22036 17464 22052
rect 17526 24028 17560 24044
rect 17526 22036 17560 22052
rect 17622 24028 17656 24044
rect 17622 22036 17656 22052
rect 16694 21968 16710 22002
rect 16744 21968 16760 22002
rect 16886 21968 16902 22002
rect 16936 21968 16952 22002
rect 17078 21968 17094 22002
rect 17128 21968 17144 22002
rect 17270 21968 17286 22002
rect 17320 21968 17336 22002
rect 17462 21968 17478 22002
rect 17512 21968 17528 22002
rect 16548 21900 16582 21962
rect 17736 21900 17770 21962
rect 16548 21866 16644 21900
rect 17674 21866 17770 21900
rect 16266 21740 17635 21775
rect 16266 21590 17370 21740
rect 17510 21590 17635 21740
rect 16266 21565 17635 21590
rect 16232 21040 16266 21102
rect 15716 21006 15812 21040
rect 16170 21006 16266 21040
rect 16656 21446 16752 21480
rect 16890 21446 16986 21480
rect 16656 21384 16690 21446
rect 14716 20586 14812 20620
rect 15554 20586 15650 20620
rect 14716 20524 14750 20586
rect 13182 19826 13278 19860
rect 14348 19826 14444 19860
rect 13182 19764 13216 19826
rect 14410 19764 14444 19826
rect 13182 16794 13216 16856
rect 15616 20524 15650 20586
rect 14958 20484 14974 20518
rect 15008 20484 15024 20518
rect 15150 20484 15166 20518
rect 15200 20484 15216 20518
rect 15342 20484 15358 20518
rect 15392 20484 15408 20518
rect 14830 20434 14864 20450
rect 14750 19172 14830 19300
rect 14926 20434 14960 20450
rect 14864 19172 14870 19300
rect 14750 19170 14870 19172
rect 14830 19156 14864 19170
rect 14926 19156 14960 19172
rect 15022 20434 15056 20450
rect 15022 19156 15056 19172
rect 15118 20434 15152 20450
rect 15118 19156 15152 19172
rect 15214 20434 15248 20450
rect 15214 19156 15248 19172
rect 15310 20434 15344 20450
rect 15310 19156 15344 19172
rect 15406 20434 15440 20450
rect 15406 19156 15440 19172
rect 15502 20434 15536 20450
rect 15502 19156 15536 19172
rect 14862 19088 14878 19122
rect 14912 19088 14928 19122
rect 15054 19088 15070 19122
rect 15104 19088 15120 19122
rect 15246 19088 15262 19122
rect 15296 19088 15312 19122
rect 15438 19088 15454 19122
rect 15488 19088 15504 19122
rect 14716 19020 14750 19082
rect 15616 19020 15650 19082
rect 14716 18986 14812 19020
rect 15554 18986 15650 19020
rect 15876 20100 15972 20134
rect 16330 20100 16426 20134
rect 15876 20038 15910 20100
rect 16392 20038 16426 20100
rect 16118 19998 16134 20032
rect 16168 19998 16184 20032
rect 15990 19948 16024 19964
rect 15990 19156 16024 19172
rect 16086 19948 16120 19964
rect 16086 19156 16120 19172
rect 16182 19948 16216 19964
rect 16182 19156 16216 19172
rect 16278 19948 16312 19964
rect 16278 19156 16312 19172
rect 16022 19088 16038 19122
rect 16072 19088 16088 19122
rect 16214 19088 16230 19122
rect 16264 19088 16280 19122
rect 15876 19020 15910 19082
rect 16392 19020 16426 19082
rect 15876 18986 15972 19020
rect 16330 18986 16426 19020
rect 16952 21384 16986 21446
rect 16656 18790 16690 18852
rect 16952 18790 16986 18852
rect 16656 18756 16752 18790
rect 16890 18756 16986 18790
rect 17020 19260 17230 21565
rect 17020 19170 17040 19260
rect 17210 19170 17230 19260
rect 14902 18634 14998 18668
rect 15156 18634 15252 18668
rect 14902 18572 14936 18634
rect 14410 16794 14444 16856
rect 13182 16760 13278 16794
rect 14348 16760 14444 16794
rect 14512 17950 14608 17984
rect 14746 17950 14842 17984
rect 14512 17888 14546 17950
rect 14808 17888 14842 17950
rect 14512 16794 14546 16856
rect 14808 16794 14842 16856
rect 14512 16760 14608 16794
rect 14746 16760 14842 16794
rect 15218 18572 15252 18634
rect 15044 18532 15060 18566
rect 15094 18532 15110 18566
rect 15016 18482 15050 18498
rect 15016 16930 15050 16946
rect 15104 18482 15138 18498
rect 15104 16930 15138 16946
rect 15044 16862 15060 16896
rect 15094 16862 15110 16896
rect 14902 16794 14936 16856
rect 15312 18634 15408 18668
rect 15566 18634 15662 18668
rect 15312 18572 15346 18634
rect 15308 18077 15312 18329
rect 15218 16794 15252 16856
rect 14902 16760 14998 16794
rect 15156 16760 15252 16794
rect 15628 18572 15662 18634
rect 15454 18532 15470 18566
rect 15504 18532 15520 18566
rect 15426 18482 15460 18498
rect 15346 18077 15426 18329
rect 15426 16930 15460 16946
rect 15514 18482 15548 18498
rect 15514 16930 15548 16946
rect 15454 16862 15470 16896
rect 15504 16862 15520 16896
rect 15312 16794 15346 16856
rect 16124 18651 16220 18685
rect 16358 18651 16454 18685
rect 16124 18589 16158 18651
rect 15628 16794 15662 16856
rect 15312 16760 15408 16794
rect 15566 16760 15662 16794
rect 15732 17950 15828 17984
rect 15966 17950 16062 17984
rect 15732 17888 15766 17950
rect 16028 17888 16062 17950
rect 15732 16794 15766 16856
rect 16028 16794 16062 16856
rect 15732 16760 15828 16794
rect 15966 16760 16062 16794
rect 16420 18589 16454 18651
rect 16124 16795 16158 16857
rect 16750 18460 16910 18756
rect 16686 18426 16782 18460
rect 16884 18426 16980 18460
rect 16686 18364 16720 18426
rect 16946 18364 16980 18426
rect 16784 18280 16800 18346
rect 16866 18280 16882 18346
rect 16686 18200 16720 18262
rect 16946 18200 16980 18262
rect 16686 18166 16782 18200
rect 16884 18166 16980 18200
rect 16420 16795 16454 16857
rect 16124 16761 16220 16795
rect 16358 16761 16454 16795
rect 17020 17280 17230 19170
rect 17266 21466 17362 21500
rect 17500 21466 17596 21500
rect 17266 21404 17300 21466
rect 17562 21404 17596 21466
rect 17266 17410 17300 17472
rect 17562 17410 17596 17472
rect 17266 17376 17362 17410
rect 17500 17376 17596 17410
rect 17020 16460 17240 17280
rect 13306 16434 17240 16460
rect 13306 16324 13326 16434
rect 13456 16334 14616 16434
rect 14736 16334 15836 16434
rect 15946 16334 17240 16434
rect 13456 16324 17240 16334
rect 13306 16308 17240 16324
rect 16941 16245 17240 16308
rect 16941 16140 17561 16245
rect 16940 16126 17561 16140
rect 14308 16044 14404 16078
rect 15242 16044 15338 16078
rect 14308 15982 14342 16044
rect 13458 15604 13554 15638
rect 13712 15604 13808 15638
rect 13458 15542 13492 15604
rect 13774 15542 13808 15604
rect 13600 15502 13616 15536
rect 13650 15502 13666 15536
rect 13572 15452 13606 15468
rect 13660 15463 13694 15468
rect 13659 15452 13774 15463
rect 13659 15327 13660 15452
rect 13572 13900 13606 13916
rect 13694 15327 13774 15452
rect 13660 13900 13694 13916
rect 13600 13832 13616 13866
rect 13650 13832 13666 13866
rect 13458 13764 13492 13826
rect 13774 13764 13808 13826
rect 13458 13730 13554 13764
rect 13712 13730 13808 13764
rect 15304 15982 15338 16044
rect 14550 15942 14566 15976
rect 14600 15942 14616 15976
rect 14742 15942 14758 15976
rect 14792 15942 14808 15976
rect 14934 15942 14950 15976
rect 14984 15942 15000 15976
rect 15126 15942 15142 15976
rect 15176 15942 15192 15976
rect 14422 15892 14456 15908
rect 14422 13900 14456 13916
rect 14518 15892 14552 15908
rect 14518 13900 14552 13916
rect 14614 15892 14648 15908
rect 14614 13900 14648 13916
rect 14710 15892 14744 15908
rect 14710 13900 14744 13916
rect 14806 15892 14840 15908
rect 14806 13900 14840 13916
rect 14902 15892 14936 15908
rect 14902 13900 14936 13916
rect 14998 15892 15032 15908
rect 14998 13900 15032 13916
rect 15094 15892 15128 15908
rect 15094 13900 15128 13916
rect 15190 15892 15224 15908
rect 15190 13900 15224 13916
rect 14454 13832 14470 13866
rect 14504 13832 14520 13866
rect 14646 13832 14662 13866
rect 14696 13832 14712 13866
rect 14838 13832 14854 13866
rect 14888 13832 14904 13866
rect 15030 13832 15046 13866
rect 15080 13832 15096 13866
rect 14308 13764 14342 13826
rect 15304 13764 15338 13826
rect 14308 13730 14404 13764
rect 15242 13730 15338 13764
rect 16018 16060 16114 16094
rect 16252 16060 16348 16094
rect 16940 16092 17074 16126
rect 17432 16093 17561 16126
rect 17432 16092 17528 16093
rect 16940 16060 17240 16092
rect 16018 15998 16052 16060
rect 16314 15998 16348 16060
rect 16018 13764 16052 13826
rect 16314 13764 16348 13826
rect 16018 13730 16114 13764
rect 16252 13730 16348 13764
rect 16978 16030 17012 16060
rect 17494 16030 17528 16092
rect 17220 15990 17236 16024
rect 17270 15990 17286 16024
rect 17092 15931 17126 15947
rect 17092 13939 17126 13955
rect 17188 15931 17222 15947
rect 17188 13939 17222 13955
rect 17284 15931 17318 15947
rect 17380 15943 17414 15947
rect 17378 15931 17494 15943
rect 17378 15824 17380 15931
rect 17284 13939 17318 13955
rect 17414 15824 17494 15931
rect 17380 13939 17414 13955
rect 17124 13862 17140 13896
rect 17174 13862 17190 13896
rect 17316 13862 17332 13896
rect 17366 13862 17382 13896
rect 16978 13794 17012 13856
rect 17528 15824 17530 15943
rect 17494 13794 17528 13856
rect 16978 13760 17074 13794
rect 17432 13760 17528 13794
rect 13074 13571 17870 13590
rect 13074 13488 13313 13571
rect 17596 13488 17870 13571
rect 13074 13455 17870 13488
rect 13074 13424 13209 13455
rect 13074 10790 13103 13424
rect 13176 10790 13209 13424
rect 17728 13433 17870 13455
rect 16122 13344 16242 13354
rect 16122 13284 16132 13344
rect 16232 13284 16242 13344
rect 13480 13195 13571 13215
rect 16122 13198 16242 13284
rect 17000 13313 17118 13334
rect 17000 13273 17021 13313
rect 17093 13273 17118 13313
rect 17000 13254 17118 13273
rect 13480 13133 13500 13195
rect 13552 13133 13571 13195
rect 13480 13115 13571 13133
rect 13614 13177 17474 13198
rect 13614 13131 13689 13177
rect 13736 13173 17474 13177
rect 13736 13131 14043 13173
rect 13614 13127 14043 13131
rect 14090 13172 15454 13173
rect 14090 13171 14749 13172
rect 14090 13127 14396 13171
rect 13614 13125 14396 13127
rect 14443 13126 14749 13171
rect 14796 13126 15100 13172
rect 15147 13127 15454 13172
rect 15501 13172 17474 13173
rect 15501 13127 15804 13172
rect 15147 13126 15804 13127
rect 15851 13171 17474 13172
rect 15851 13126 16156 13171
rect 14443 13125 16156 13126
rect 16203 13125 16509 13171
rect 16556 13125 16858 13171
rect 16905 13125 17212 13171
rect 17259 13125 17385 13171
rect 17432 13125 17474 13171
rect 13614 13119 17474 13125
rect 13675 13115 13750 13119
rect 14029 13111 14104 13119
rect 14382 13109 14457 13119
rect 14735 13110 14810 13119
rect 15086 13110 15161 13119
rect 15440 13111 15515 13119
rect 15790 13110 15865 13119
rect 16122 13114 16242 13119
rect 16142 13109 16217 13114
rect 16495 13109 16570 13119
rect 16844 13109 16919 13119
rect 17198 13109 17273 13119
rect 17371 13109 17446 13119
rect 13434 13058 13468 13074
rect 13434 11066 13468 11082
rect 13522 13058 13556 13074
rect 13522 11066 13556 11082
rect 13610 13058 13644 13074
rect 13610 11066 13644 11082
rect 13698 13058 13732 13074
rect 13698 11066 13732 11082
rect 13786 13058 13820 13074
rect 13786 11066 13820 11082
rect 13874 13058 13908 13074
rect 13874 11066 13908 11082
rect 13962 13058 13996 13074
rect 13962 11066 13996 11082
rect 14050 13058 14084 13074
rect 14050 11066 14084 11082
rect 14138 13058 14172 13074
rect 14138 11066 14172 11082
rect 14226 13058 14260 13074
rect 14226 11066 14260 11082
rect 14314 13058 14348 13074
rect 14314 11066 14348 11082
rect 14402 13058 14436 13074
rect 14402 11066 14436 11082
rect 14490 13058 14524 13074
rect 14490 11066 14524 11082
rect 14578 13058 14612 13074
rect 14578 11066 14612 11082
rect 14666 13058 14700 13074
rect 14666 11066 14700 11082
rect 14754 13058 14788 13074
rect 14754 11066 14788 11082
rect 14842 13058 14876 13074
rect 14842 11066 14876 11082
rect 14930 13058 14964 13074
rect 14930 11066 14964 11082
rect 15018 13058 15052 13074
rect 15018 11066 15052 11082
rect 15106 13058 15140 13074
rect 15106 11066 15140 11082
rect 15194 13058 15228 13074
rect 15194 11066 15228 11082
rect 15282 13058 15316 13074
rect 15282 11066 15316 11082
rect 15370 13058 15404 13074
rect 15370 11066 15404 11082
rect 15458 13058 15492 13074
rect 15458 11066 15492 11082
rect 15546 13058 15580 13074
rect 15546 11066 15580 11082
rect 15634 13058 15668 13074
rect 15634 11066 15668 11082
rect 15722 13058 15756 13074
rect 15722 11066 15756 11082
rect 15810 13058 15844 13074
rect 15810 11066 15844 11082
rect 15898 13058 15932 13074
rect 15898 11066 15932 11082
rect 15986 13058 16020 13074
rect 15986 11066 16020 11082
rect 16074 13058 16108 13074
rect 16074 11066 16108 11082
rect 16162 13058 16196 13074
rect 16162 11066 16196 11082
rect 16250 13058 16284 13074
rect 16250 11066 16284 11082
rect 16338 13058 16372 13074
rect 16338 11066 16372 11082
rect 16426 13058 16460 13074
rect 16426 11066 16460 11082
rect 16514 13058 16548 13074
rect 16514 11066 16548 11082
rect 16602 13058 16636 13074
rect 16602 11066 16636 11082
rect 16690 13058 16724 13074
rect 16690 11066 16724 11082
rect 16778 13058 16812 13074
rect 16778 11066 16812 11082
rect 16866 13058 16900 13074
rect 16866 11066 16900 11082
rect 16954 13058 16988 13074
rect 16954 11066 16988 11082
rect 17042 13058 17076 13074
rect 17042 11066 17076 11082
rect 17130 13058 17164 13074
rect 17130 11066 17164 11082
rect 17218 13058 17252 13074
rect 17218 11066 17252 11082
rect 17306 13058 17340 13074
rect 17306 11066 17340 11082
rect 17394 13058 17428 13074
rect 17394 11066 17428 11082
rect 17482 13058 17516 13074
rect 17482 11066 17516 11082
rect 13497 11002 13572 11020
rect 13497 11000 13511 11002
rect 13467 10956 13511 11000
rect 13558 11000 13572 11002
rect 13847 11000 13922 11014
rect 14205 11000 14280 11017
rect 14553 11000 14628 11017
rect 14904 11000 14979 11017
rect 15255 11000 15330 11016
rect 15606 11000 15681 11014
rect 15961 11000 16036 11017
rect 16311 11000 16386 11013
rect 16665 11000 16740 11015
rect 17015 11000 17090 11013
rect 13558 10999 17158 11000
rect 13558 10996 14219 10999
rect 13558 10956 13861 10996
rect 13467 10950 13861 10956
rect 13908 10953 14219 10996
rect 14266 10953 14567 10999
rect 14614 10953 14918 10999
rect 14965 10998 15975 10999
rect 14965 10953 15269 10998
rect 13908 10952 15269 10953
rect 15316 10996 15975 10998
rect 15316 10952 15620 10996
rect 13908 10950 15620 10952
rect 15667 10953 15975 10996
rect 16022 10997 17158 10999
rect 16022 10995 16679 10997
rect 16022 10953 16325 10995
rect 15667 10950 16325 10953
rect 13467 10949 16325 10950
rect 16372 10951 16679 10995
rect 16726 10995 17158 10997
rect 16726 10951 17029 10995
rect 16372 10949 17029 10951
rect 17076 10949 17158 10995
rect 13467 10931 17158 10949
rect 17352 10994 17472 11024
rect 13467 10874 13597 10931
rect 17352 10914 17372 10994
rect 17452 10914 17472 10994
rect 17352 10894 17472 10914
rect 13467 10815 13482 10874
rect 13581 10815 13597 10874
rect 13467 10804 13597 10815
rect 17342 10874 17482 10894
rect 13074 10738 13209 10790
rect 17342 10784 17362 10874
rect 17462 10784 17482 10874
rect 17342 10774 17482 10784
rect 17728 10799 17766 13433
rect 17839 10799 17870 13433
rect 17728 10738 17870 10799
rect 13074 10718 17870 10738
rect 13074 10635 13355 10718
rect 17638 10635 17870 10718
rect 13074 10610 17870 10635
rect 13861 10532 17005 10610
rect 13850 9688 17008 10532
rect 13850 8938 13906 9688
rect 16938 8938 17008 9688
rect 13850 8882 17008 8938
<< viali >>
rect 14118 27684 16404 28832
rect 13064 24562 13461 24600
rect 16495 24562 16892 24600
rect 13094 23882 13491 23920
rect 14325 23882 14722 23920
rect 13090 23390 13310 23550
rect 16290 23430 16430 23560
rect 13502 21655 13540 22052
rect 13502 21124 13540 21521
rect 14114 23188 14148 23222
rect 14306 23188 14340 23222
rect 14498 23188 14532 23222
rect 14690 23188 14724 23222
rect 13970 21162 14004 23138
rect 14066 21162 14100 23138
rect 14162 21162 14196 23138
rect 14258 21162 14292 23138
rect 14354 21162 14388 23138
rect 14450 21162 14484 23138
rect 14546 21162 14580 23138
rect 14642 21162 14676 23138
rect 14738 21162 14772 23138
rect 14830 23040 14852 23140
rect 14852 23040 14886 23140
rect 14886 23040 14900 23140
rect 14018 21078 14052 21112
rect 14210 21078 14244 21112
rect 14402 21078 14436 21112
rect 14594 21078 14628 21112
rect 15322 22815 15360 23212
rect 15322 21144 15360 21541
rect 15974 23236 16008 23270
rect 15830 21201 15864 23177
rect 15926 21201 15960 23177
rect 16022 21201 16056 23177
rect 16118 21201 16152 23177
rect 15878 21108 15912 21142
rect 16070 21108 16104 21142
rect 16806 24078 16840 24112
rect 16998 24078 17032 24112
rect 17190 24078 17224 24112
rect 17382 24078 17416 24112
rect 17574 24078 17608 24112
rect 16662 22052 16696 24028
rect 16758 22052 16792 24028
rect 16854 22052 16888 24028
rect 16950 22052 16984 24028
rect 17046 22052 17080 24028
rect 17142 22052 17176 24028
rect 17238 22052 17272 24028
rect 17334 22052 17368 24028
rect 17430 22052 17464 24028
rect 17526 22052 17560 24028
rect 17622 22052 17656 24028
rect 16710 21968 16744 22002
rect 16902 21968 16936 22002
rect 17094 21968 17128 22002
rect 17286 21968 17320 22002
rect 17478 21968 17512 22002
rect 17370 21590 17510 21740
rect 13330 19608 13727 19714
rect 13899 19608 14296 19714
rect 13330 19222 13727 19328
rect 13899 19222 14296 19328
rect 13330 18836 13727 18942
rect 13899 18836 14296 18942
rect 13330 18450 13727 18556
rect 13899 18450 14296 18556
rect 13330 18064 13727 18170
rect 13899 18064 14296 18170
rect 13330 17678 13727 17784
rect 13899 17678 14296 17784
rect 13330 17292 13727 17398
rect 13899 17292 14296 17398
rect 13330 16906 13727 17012
rect 13899 16906 14296 17012
rect 14974 20484 15008 20518
rect 15166 20484 15200 20518
rect 15358 20484 15392 20518
rect 14830 19172 14864 20434
rect 14926 19172 14960 20434
rect 15022 19172 15056 20434
rect 15118 19172 15152 20434
rect 15214 19172 15248 20434
rect 15310 19172 15344 20434
rect 15406 19172 15440 20434
rect 15502 19172 15536 20434
rect 14878 19088 14912 19122
rect 15070 19088 15104 19122
rect 15262 19088 15296 19122
rect 15454 19088 15488 19122
rect 16134 19998 16168 20032
rect 15990 19172 16024 19948
rect 16086 19172 16120 19948
rect 16182 19172 16216 19948
rect 16278 19172 16312 19948
rect 16038 19088 16072 19122
rect 16230 19088 16264 19122
rect 16802 20935 16840 21332
rect 16802 18904 16840 19301
rect 17040 19170 17210 19260
rect 14658 17439 14696 17836
rect 14658 16908 14696 17305
rect 15060 18532 15094 18566
rect 15016 16946 15050 18482
rect 15104 16946 15138 18482
rect 15060 16862 15094 16896
rect 15470 18532 15504 18566
rect 15426 16946 15460 18482
rect 15514 16946 15548 18482
rect 15470 16862 15504 16896
rect 15878 17439 15916 17836
rect 15878 16908 15916 17305
rect 16270 18140 16308 18537
rect 16270 16909 16308 17306
rect 16800 18280 16866 18346
rect 17412 20955 17450 21352
rect 17412 17524 17450 17921
rect 13326 16324 13456 16434
rect 14616 16334 14736 16434
rect 15836 16334 15946 16434
rect 13616 15502 13650 15536
rect 13572 13916 13606 15452
rect 13660 13916 13694 15452
rect 13616 13832 13650 13866
rect 14566 15942 14600 15976
rect 14758 15942 14792 15976
rect 14950 15942 14984 15976
rect 15142 15942 15176 15976
rect 14422 13916 14456 15892
rect 14518 13916 14552 15892
rect 14614 13916 14648 15892
rect 14710 13916 14744 15892
rect 14806 13916 14840 15892
rect 14902 13916 14936 15892
rect 14998 13916 15032 15892
rect 15094 13916 15128 15892
rect 15190 13916 15224 15892
rect 14470 13832 14504 13866
rect 14662 13832 14696 13866
rect 14854 13832 14888 13866
rect 15046 13832 15080 13866
rect 16164 15549 16202 15946
rect 16164 13878 16202 14275
rect 17236 15990 17270 16024
rect 17092 13955 17126 15931
rect 17188 13955 17222 15931
rect 17284 13955 17318 15931
rect 17380 13955 17414 15931
rect 17140 13862 17174 13896
rect 17332 13862 17366 13896
rect 16132 13284 16232 13344
rect 17021 13273 17093 13313
rect 13500 13133 13552 13195
rect 13434 11082 13468 13058
rect 13522 11082 13556 13058
rect 13610 11082 13644 13058
rect 13698 11082 13732 13058
rect 13786 11082 13820 13058
rect 13874 11082 13908 13058
rect 13962 11082 13996 13058
rect 14050 11082 14084 13058
rect 14138 11082 14172 13058
rect 14226 11082 14260 13058
rect 14314 11082 14348 13058
rect 14402 11082 14436 13058
rect 14490 11082 14524 13058
rect 14578 11082 14612 13058
rect 14666 11082 14700 13058
rect 14754 11082 14788 13058
rect 14842 11082 14876 13058
rect 14930 11082 14964 13058
rect 15018 11082 15052 13058
rect 15106 11082 15140 13058
rect 15194 11082 15228 13058
rect 15282 11082 15316 13058
rect 15370 11082 15404 13058
rect 15458 11082 15492 13058
rect 15546 11082 15580 13058
rect 15634 11082 15668 13058
rect 15722 11082 15756 13058
rect 15810 11082 15844 13058
rect 15898 11082 15932 13058
rect 15986 11082 16020 13058
rect 16074 11082 16108 13058
rect 16162 11082 16196 13058
rect 16250 11082 16284 13058
rect 16338 11082 16372 13058
rect 16426 11082 16460 13058
rect 16514 11082 16548 13058
rect 16602 11082 16636 13058
rect 16690 11082 16724 13058
rect 16778 11082 16812 13058
rect 16866 11082 16900 13058
rect 16954 11082 16988 13058
rect 17042 11082 17076 13058
rect 17130 11082 17164 13058
rect 17218 11082 17252 13058
rect 17306 11082 17340 13058
rect 17394 11082 17428 13058
rect 17482 11082 17516 13058
rect 13482 10815 13581 10874
rect 17362 10784 17462 10874
rect 14502 10654 14682 10714
rect 13906 8938 16938 9688
<< metal1 >>
rect 2229 28892 28685 28930
rect 2229 28832 27180 28892
rect 2229 28820 14118 28832
rect 2229 27686 2340 28820
rect 3694 27686 14118 28820
rect 2229 27684 14118 27686
rect 16404 27758 27180 28832
rect 28534 27758 28685 28892
rect 16404 27684 28685 27758
rect 2229 27600 28685 27684
rect 4162 26962 26614 26978
rect 4162 26954 25304 26962
rect 4162 25634 4246 26954
rect 5518 25642 25304 26954
rect 26576 25642 26614 26962
rect 5518 25634 26614 25642
rect 4162 25554 26614 25634
rect 16810 24610 16910 24620
rect 16810 24606 16820 24610
rect 13052 24600 13473 24606
rect 13052 24562 13064 24600
rect 13461 24562 13473 24600
rect 13052 24556 13473 24562
rect 16483 24600 16820 24606
rect 16483 24562 16495 24600
rect 16483 24556 16820 24562
rect 16810 24520 16820 24556
rect 16900 24520 16910 24610
rect 16810 24510 16910 24520
rect 12535 24142 16435 24280
rect 12535 24140 16441 24142
rect 12535 24112 17620 24140
rect 12535 24078 16806 24112
rect 16840 24078 16998 24112
rect 17032 24078 17190 24112
rect 17224 24078 17382 24112
rect 17416 24078 17574 24112
rect 17608 24078 17620 24112
rect 12535 24070 17620 24078
rect 12535 24003 16441 24070
rect 12535 17968 12812 24003
rect 13070 23926 13340 23940
rect 13070 23920 13503 23926
rect 13070 23882 13094 23920
rect 13491 23882 13503 23920
rect 13070 23876 13503 23882
rect 14303 23920 16441 24003
rect 14303 23882 14325 23920
rect 14722 23882 16441 23920
rect 13070 23550 13340 23876
rect 14303 23865 16441 23882
rect 16656 24028 16702 24040
rect 13070 23390 13090 23550
rect 13310 23390 13340 23550
rect 13070 23370 13340 23390
rect 15260 23612 15432 23632
rect 13648 23372 13802 23388
rect 13648 23042 13664 23372
rect 13792 23042 13802 23372
rect 15260 23364 15272 23612
rect 15414 23364 15432 23612
rect 16270 23560 16450 23580
rect 16270 23430 16290 23560
rect 16430 23430 16450 23560
rect 16270 23410 16450 23430
rect 15260 23312 15432 23364
rect 14090 23222 14740 23240
rect 14090 23188 14114 23222
rect 14148 23188 14306 23222
rect 14340 23188 14498 23222
rect 14532 23188 14690 23222
rect 14724 23188 14740 23222
rect 14090 23180 14740 23188
rect 15260 23212 15420 23312
rect 15950 23270 16030 23280
rect 15950 23236 15974 23270
rect 16008 23236 16030 23270
rect 15950 23230 16030 23236
rect 13648 23028 13802 23042
rect 13964 23138 14010 23150
rect 13496 22052 13546 22064
rect 13496 21780 13502 22052
rect 13480 21655 13502 21780
rect 13540 21780 13546 22052
rect 13650 21780 13800 23028
rect 13540 21655 13800 21780
rect 13480 21630 13800 21655
rect 13496 21521 13546 21533
rect 13496 21190 13502 21521
rect 12535 17700 12559 17968
rect 12791 17700 12812 17968
rect 12535 17676 12812 17700
rect 13000 21124 13502 21190
rect 13540 21190 13546 21521
rect 13540 21124 13560 21190
rect 13000 21070 13560 21124
rect 13710 21120 13800 21630
rect 13964 21271 13970 23138
rect 13951 21252 13970 21271
rect 14004 21271 14010 23138
rect 14041 23138 14111 23151
rect 14041 23132 14066 23138
rect 14100 23132 14111 23138
rect 14041 23050 14050 23132
rect 14102 23050 14111 23132
rect 14041 23031 14066 23050
rect 14004 21252 14021 21271
rect 13951 21170 13960 21252
rect 14012 21170 14021 21252
rect 13951 21162 13970 21170
rect 14004 21162 14021 21170
rect 13951 21151 14021 21162
rect 14060 21162 14066 23031
rect 14100 23031 14111 23050
rect 14156 23138 14202 23150
rect 14100 21162 14106 23031
rect 14156 21271 14162 23138
rect 13964 21150 14010 21151
rect 14060 21150 14106 21162
rect 14141 21252 14162 21271
rect 14196 21271 14202 23138
rect 14241 23138 14311 23151
rect 14241 23132 14258 23138
rect 14292 23132 14311 23138
rect 14241 23050 14250 23132
rect 14302 23050 14311 23132
rect 14241 23031 14258 23050
rect 14196 21252 14211 21271
rect 14141 21170 14150 21252
rect 14202 21170 14211 21252
rect 14141 21162 14162 21170
rect 14196 21162 14211 21170
rect 14141 21151 14211 21162
rect 14252 21162 14258 23031
rect 14292 23031 14311 23050
rect 14348 23138 14394 23150
rect 14292 21162 14298 23031
rect 14348 21271 14354 23138
rect 14156 21150 14202 21151
rect 14252 21150 14298 21162
rect 14331 21252 14354 21271
rect 14388 21271 14394 23138
rect 14431 23138 14501 23151
rect 14431 23132 14450 23138
rect 14484 23132 14501 23138
rect 14431 23050 14440 23132
rect 14492 23050 14501 23132
rect 14431 23031 14450 23050
rect 14388 21252 14401 21271
rect 14331 21170 14340 21252
rect 14392 21170 14401 21252
rect 14331 21162 14354 21170
rect 14388 21162 14401 21170
rect 14331 21151 14401 21162
rect 14444 21162 14450 23031
rect 14484 23031 14501 23050
rect 14540 23138 14586 23150
rect 14484 21162 14490 23031
rect 14540 21271 14546 23138
rect 14348 21150 14394 21151
rect 14444 21150 14490 21162
rect 14521 21252 14546 21271
rect 14580 21271 14586 23138
rect 14621 23138 14691 23151
rect 14621 23132 14642 23138
rect 14676 23132 14691 23138
rect 14621 23050 14630 23132
rect 14682 23050 14691 23132
rect 14621 23031 14642 23050
rect 14580 21252 14591 21271
rect 14521 21170 14530 21252
rect 14582 21170 14591 21252
rect 14521 21162 14546 21170
rect 14580 21162 14591 21170
rect 14521 21151 14591 21162
rect 14636 21162 14642 23031
rect 14676 23031 14691 23050
rect 14732 23138 14778 23150
rect 14676 21162 14682 23031
rect 14732 21271 14738 23138
rect 14540 21150 14586 21151
rect 14636 21150 14682 21162
rect 14721 21252 14738 21271
rect 14772 21271 14778 23138
rect 14810 23140 14920 23160
rect 14810 23040 14830 23140
rect 14900 23040 14920 23140
rect 14810 23020 14920 23040
rect 15260 22815 15322 23212
rect 15360 22815 15420 23212
rect 15260 22760 15420 22815
rect 15824 23177 15870 23189
rect 15316 21541 15366 21553
rect 15316 21290 15322 21541
rect 14772 21252 14791 21271
rect 14721 21170 14730 21252
rect 14782 21170 14791 21252
rect 14721 21162 14738 21170
rect 14772 21162 14791 21170
rect 14721 21151 14791 21162
rect 14732 21150 14778 21151
rect 15290 21144 15322 21290
rect 15360 21290 15366 21541
rect 15824 21311 15830 23177
rect 15801 21292 15830 21311
rect 15864 21311 15870 23177
rect 15901 23177 15971 23191
rect 15901 23172 15926 23177
rect 15960 23172 15971 23177
rect 15901 23090 15910 23172
rect 15962 23090 15971 23172
rect 15901 23071 15926 23090
rect 15360 21150 15390 21290
rect 15801 21210 15810 21292
rect 15801 21201 15830 21210
rect 15864 21201 15871 21311
rect 15801 21191 15871 21201
rect 15920 21201 15926 23071
rect 15960 23071 15971 23090
rect 16016 23177 16062 23189
rect 15960 21201 15966 23071
rect 16016 21311 16022 23177
rect 15824 21189 15870 21191
rect 15920 21189 15966 21201
rect 16001 21292 16022 21311
rect 16056 21311 16062 23177
rect 16091 23177 16161 23191
rect 16091 23172 16118 23177
rect 16091 23090 16100 23172
rect 16091 23071 16118 23090
rect 16056 21292 16071 21311
rect 16001 21210 16010 21292
rect 16062 21210 16071 21292
rect 16001 21201 16022 21210
rect 16056 21201 16071 21210
rect 16001 21191 16071 21201
rect 16112 21201 16118 23071
rect 16152 23071 16161 23177
rect 16152 21201 16158 23071
rect 16656 22170 16662 24028
rect 16651 22160 16662 22170
rect 16696 22170 16702 24028
rect 16743 24031 16813 24041
rect 16743 23920 16750 24031
rect 16803 23920 16813 24031
rect 16743 23911 16758 23920
rect 16696 22160 16721 22170
rect 16651 22049 16658 22160
rect 16711 22049 16721 22160
rect 16651 22040 16721 22049
rect 16752 22052 16758 23911
rect 16792 23911 16813 23920
rect 16848 24028 16894 24040
rect 16792 22052 16798 23911
rect 16848 22170 16854 24028
rect 16752 22040 16798 22052
rect 16832 22160 16854 22170
rect 16888 22170 16894 24028
rect 16933 24031 17003 24041
rect 16933 23920 16940 24031
rect 16993 23920 17003 24031
rect 16933 23911 16950 23920
rect 16888 22160 16902 22170
rect 16832 22049 16839 22160
rect 16892 22049 16902 22160
rect 16832 22040 16902 22049
rect 16944 22052 16950 23911
rect 16984 23911 17003 23920
rect 17040 24028 17086 24040
rect 16984 22052 16990 23911
rect 17040 22170 17046 24028
rect 16944 22040 16990 22052
rect 17022 22160 17046 22170
rect 17080 22170 17086 24028
rect 17123 24031 17193 24041
rect 17123 23920 17130 24031
rect 17183 23920 17193 24031
rect 17123 23911 17142 23920
rect 17080 22160 17092 22170
rect 17022 22049 17029 22160
rect 17082 22049 17092 22160
rect 17022 22040 17092 22049
rect 17136 22052 17142 23911
rect 17176 23911 17193 23920
rect 17232 24028 17278 24040
rect 17176 22052 17182 23911
rect 17232 22173 17238 24028
rect 17136 22040 17182 22052
rect 17213 22163 17238 22173
rect 17272 22173 17278 24028
rect 17313 24031 17383 24041
rect 17313 23920 17320 24031
rect 17373 23920 17383 24031
rect 17313 23911 17334 23920
rect 17272 22163 17283 22173
rect 17213 22052 17220 22163
rect 17273 22052 17283 22163
rect 17213 22043 17283 22052
rect 17328 22052 17334 23911
rect 17368 23911 17383 23920
rect 17424 24028 17470 24040
rect 17368 22052 17374 23911
rect 17424 22171 17430 24028
rect 17232 22040 17278 22043
rect 17328 22040 17374 22052
rect 17412 22161 17430 22171
rect 17464 22171 17470 24028
rect 17513 24031 17583 24041
rect 17513 23920 17520 24031
rect 17573 23920 17583 24031
rect 17513 23911 17526 23920
rect 17464 22161 17482 22171
rect 17412 22050 17419 22161
rect 17472 22050 17482 22161
rect 17412 22041 17482 22050
rect 17520 22052 17526 23911
rect 17560 23911 17583 23920
rect 17616 24028 17662 24040
rect 17560 22052 17566 23911
rect 17616 22172 17622 24028
rect 17424 22040 17470 22041
rect 17520 22040 17566 22052
rect 17603 22162 17622 22172
rect 17656 22172 17662 24028
rect 17656 22162 17673 22172
rect 17603 22051 17610 22162
rect 17663 22051 17673 22162
rect 17603 22042 17673 22051
rect 17616 22040 17662 22042
rect 16690 22002 17530 22010
rect 16690 21968 16710 22002
rect 16744 21968 16902 22002
rect 16936 21968 17094 22002
rect 17128 21968 17286 22002
rect 17320 21968 17478 22002
rect 17512 21968 17530 22002
rect 16690 21940 17530 21968
rect 17350 21740 17530 21770
rect 17350 21590 17370 21740
rect 17510 21590 17530 21740
rect 17350 21370 17530 21590
rect 17390 21352 17480 21370
rect 16016 21189 16062 21191
rect 16112 21189 16158 21201
rect 16780 21332 17130 21350
rect 15360 21144 16120 21150
rect 15290 21142 16120 21144
rect 13710 21112 14650 21120
rect 13710 21078 14018 21112
rect 14052 21078 14210 21112
rect 14244 21078 14402 21112
rect 14436 21078 14594 21112
rect 14628 21078 14650 21112
rect 15290 21108 15878 21142
rect 15912 21108 16070 21142
rect 16104 21108 16120 21142
rect 15290 21080 16120 21108
rect 13000 16224 13120 21070
rect 13710 21040 14650 21078
rect 16780 20935 16802 21332
rect 16840 21322 17130 21332
rect 16840 20935 16864 21322
rect 16780 20932 16864 20935
rect 17006 20932 17130 21322
rect 17390 21070 17412 21352
rect 17406 20955 17412 21070
rect 17450 21070 17480 21352
rect 17450 20955 17456 21070
rect 17406 20943 17456 20955
rect 16780 20910 17130 20932
rect 14880 20550 15490 20570
rect 14880 20490 14920 20550
rect 15460 20490 15490 20550
rect 14880 20484 14974 20490
rect 15008 20484 15166 20490
rect 15200 20484 15358 20490
rect 15392 20484 15490 20490
rect 14880 20480 15490 20484
rect 14962 20478 15020 20480
rect 15154 20478 15212 20480
rect 15346 20478 15404 20480
rect 14824 20434 14870 20446
rect 14920 20440 14966 20446
rect 13306 19720 13486 19734
rect 14136 19720 14316 19734
rect 13306 19714 13739 19720
rect 13306 19608 13330 19714
rect 13727 19608 13739 19714
rect 13306 19602 13739 19608
rect 13887 19714 14316 19720
rect 13887 19608 13899 19714
rect 14296 19608 14316 19714
rect 13887 19602 14316 19608
rect 13306 19334 13486 19602
rect 14136 19334 14316 19602
rect 13306 19328 13739 19334
rect 13306 19222 13330 19328
rect 13727 19222 13739 19328
rect 13306 19216 13739 19222
rect 13887 19328 14316 19334
rect 13887 19222 13899 19328
rect 14296 19222 14316 19328
rect 14824 19300 14830 20434
rect 13887 19216 14316 19222
rect 13306 18948 13486 19216
rect 14136 18948 14316 19216
rect 14810 19290 14830 19300
rect 14864 19300 14870 20434
rect 14900 20434 14980 20440
rect 14900 20430 14926 20434
rect 14960 20430 14980 20434
rect 14900 20320 14910 20430
rect 14970 20320 14980 20430
rect 14900 20310 14926 20320
rect 14864 19290 14890 19300
rect 14810 19180 14820 19290
rect 14880 19180 14890 19290
rect 14810 19172 14830 19180
rect 14864 19172 14890 19180
rect 14810 19170 14890 19172
rect 14920 19172 14926 20310
rect 14960 20310 14980 20320
rect 15016 20434 15062 20446
rect 15112 20440 15158 20446
rect 14960 19172 14966 20310
rect 15016 19300 15022 20434
rect 14824 19160 14870 19170
rect 14920 19160 14966 19172
rect 15000 19290 15022 19300
rect 15056 19300 15062 20434
rect 15090 20434 15170 20440
rect 15090 20430 15118 20434
rect 15152 20430 15170 20434
rect 15090 20320 15100 20430
rect 15160 20320 15170 20430
rect 15090 20310 15118 20320
rect 15056 19290 15080 19300
rect 15000 19180 15010 19290
rect 15070 19180 15080 19290
rect 15000 19172 15022 19180
rect 15056 19172 15080 19180
rect 15000 19170 15080 19172
rect 15112 19172 15118 20310
rect 15152 20310 15170 20320
rect 15208 20434 15254 20446
rect 15304 20440 15350 20446
rect 15152 19172 15158 20310
rect 15208 19300 15214 20434
rect 15016 19160 15062 19170
rect 15112 19160 15158 19172
rect 15190 19290 15214 19300
rect 15248 19300 15254 20434
rect 15290 20434 15370 20440
rect 15290 20430 15310 20434
rect 15344 20430 15370 20434
rect 15290 20320 15300 20430
rect 15360 20320 15370 20430
rect 15290 20310 15310 20320
rect 15248 19290 15270 19300
rect 15190 19180 15200 19290
rect 15260 19180 15270 19290
rect 15190 19172 15214 19180
rect 15248 19172 15270 19180
rect 15190 19170 15270 19172
rect 15304 19172 15310 20310
rect 15344 20310 15370 20320
rect 15400 20434 15446 20446
rect 15496 20440 15542 20446
rect 15344 19172 15350 20310
rect 15400 19300 15406 20434
rect 15208 19160 15254 19170
rect 15304 19160 15350 19172
rect 15380 19290 15406 19300
rect 15440 19300 15446 20434
rect 15480 20434 15560 20440
rect 15480 20430 15502 20434
rect 15536 20430 15560 20434
rect 15480 20320 15490 20430
rect 15550 20320 15560 20430
rect 15480 20310 15502 20320
rect 15440 19290 15460 19300
rect 15380 19180 15390 19290
rect 15450 19180 15460 19290
rect 15380 19172 15406 19180
rect 15440 19172 15460 19180
rect 15380 19170 15460 19172
rect 15496 19172 15502 20310
rect 15536 20310 15560 20320
rect 15536 19172 15542 20310
rect 16120 20032 16180 20050
rect 16120 19998 16134 20032
rect 16168 19998 16180 20032
rect 16120 19990 16180 19998
rect 15984 19948 16030 19960
rect 15984 19290 15990 19948
rect 15400 19160 15446 19170
rect 15496 19160 15542 19172
rect 15960 19280 15990 19290
rect 16024 19290 16030 19948
rect 16060 19950 16140 19960
rect 16060 19840 16070 19950
rect 16130 19840 16140 19950
rect 16060 19830 16086 19840
rect 16024 19280 16040 19290
rect 15960 19170 15970 19280
rect 16030 19170 16040 19280
rect 15960 19160 16040 19170
rect 16080 19172 16086 19830
rect 16120 19830 16140 19840
rect 16176 19948 16222 19960
rect 16120 19172 16126 19830
rect 16176 19290 16182 19948
rect 16080 19160 16126 19172
rect 16160 19280 16182 19290
rect 16216 19290 16222 19948
rect 16250 19950 16330 19960
rect 16250 19840 16260 19950
rect 16320 19840 16330 19950
rect 16250 19830 16278 19840
rect 16216 19280 16240 19290
rect 16160 19170 16170 19280
rect 16230 19170 16240 19280
rect 16160 19160 16240 19170
rect 16272 19172 16278 19830
rect 16312 19830 16330 19840
rect 16312 19172 16318 19830
rect 16272 19160 16318 19172
rect 16796 19301 16846 19313
rect 14860 19122 15510 19130
rect 14860 19088 14878 19122
rect 14912 19088 15070 19122
rect 15104 19088 15262 19122
rect 15296 19088 15454 19122
rect 15488 19088 15510 19122
rect 14860 19060 15510 19088
rect 16020 19122 16610 19130
rect 16020 19088 16038 19122
rect 16072 19088 16230 19122
rect 16264 19120 16610 19122
rect 16264 19088 16500 19120
rect 16020 19070 16500 19088
rect 13306 18942 13739 18948
rect 13306 18836 13330 18942
rect 13727 18836 13739 18942
rect 13306 18830 13739 18836
rect 13887 18942 14316 18948
rect 13887 18836 13899 18942
rect 14296 18836 14316 18942
rect 15140 18980 15260 19060
rect 16490 19030 16500 19070
rect 16600 19030 16610 19120
rect 16490 19020 16610 19030
rect 16796 18980 16802 19301
rect 15140 18904 16802 18980
rect 16840 18980 16846 19301
rect 17020 19260 17230 19280
rect 17020 19170 17040 19260
rect 17210 19170 17230 19260
rect 17020 19160 17230 19170
rect 16840 18904 16860 18980
rect 15140 18860 16860 18904
rect 13887 18830 14316 18836
rect 13306 18562 13486 18830
rect 14136 18562 14316 18830
rect 15038 18714 16326 18787
rect 15038 18584 15111 18714
rect 13306 18556 13739 18562
rect 13306 18450 13330 18556
rect 13727 18450 13739 18556
rect 13306 18444 13739 18450
rect 13887 18556 14316 18562
rect 13887 18450 13899 18556
rect 14296 18450 14316 18556
rect 15036 18566 15116 18584
rect 15036 18532 15060 18566
rect 15094 18532 15116 18566
rect 15036 18524 15116 18532
rect 15446 18566 15526 18584
rect 15446 18532 15470 18566
rect 15504 18532 15526 18566
rect 15446 18524 15526 18532
rect 16253 18537 16326 18714
rect 13887 18444 14316 18450
rect 13306 18176 13486 18444
rect 14136 18176 14316 18444
rect 15010 18482 15056 18494
rect 15010 18209 15016 18482
rect 13306 18170 13739 18176
rect 13306 18064 13330 18170
rect 13727 18064 13739 18170
rect 13306 18058 13739 18064
rect 13887 18170 14316 18176
rect 13887 18064 13899 18170
rect 14296 18064 14316 18170
rect 13887 18058 14316 18064
rect 13306 17790 13486 18058
rect 14136 17790 14316 18058
rect 13306 17784 13739 17790
rect 13306 17678 13330 17784
rect 13727 17678 13739 17784
rect 13306 17672 13739 17678
rect 13887 17784 14316 17790
rect 13887 17678 13899 17784
rect 14296 17678 14316 17784
rect 13887 17672 14316 17678
rect 13306 17404 13486 17672
rect 14136 17404 14316 17672
rect 13306 17398 13739 17404
rect 13306 17292 13330 17398
rect 13727 17292 13739 17398
rect 13306 17286 13739 17292
rect 13887 17398 14316 17404
rect 13887 17292 13899 17398
rect 14296 17292 14316 17398
rect 13887 17286 14316 17292
rect 13306 17018 13486 17286
rect 14136 17018 14316 17286
rect 13306 17012 13739 17018
rect 13306 16906 13330 17012
rect 13727 16906 13739 17012
rect 13306 16900 13739 16906
rect 13887 17012 14316 17018
rect 13887 16906 13899 17012
rect 14296 16906 14316 17012
rect 13887 16900 14316 16906
rect 13306 16434 13486 16900
rect 14136 16694 14316 16900
rect 14136 16574 14156 16694
rect 14286 16574 14316 16694
rect 14136 16554 14316 16574
rect 14371 18096 15016 18209
rect 13306 16324 13326 16434
rect 13456 16324 13486 16434
rect 13306 16304 13486 16324
rect 13516 16392 13612 16397
rect 14371 16392 14484 18096
rect 14641 17836 14755 17851
rect 14641 17833 14658 17836
rect 14696 17833 14755 17836
rect 14641 17606 14654 17833
rect 14737 17606 14755 17833
rect 14641 17594 14658 17606
rect 14652 17439 14658 17594
rect 14696 17594 14755 17606
rect 14696 17439 14702 17594
rect 14652 17427 14702 17439
rect 14652 17305 14702 17317
rect 14652 17004 14658 17305
rect 13516 16384 14484 16392
rect 13516 16289 13528 16384
rect 13592 16289 14484 16384
rect 14596 16908 14658 17004
rect 14696 17004 14702 17305
rect 14696 16908 14756 17004
rect 15010 16946 15016 18096
rect 15050 16946 15056 18482
rect 15010 16934 15056 16946
rect 15098 18482 15144 18494
rect 15098 16946 15104 18482
rect 15138 17851 15144 18482
rect 15420 18482 15466 18494
rect 15138 17835 15187 17851
rect 15175 17606 15187 17835
rect 15138 17596 15187 17606
rect 15138 17044 15144 17596
rect 15138 16946 15265 17044
rect 15098 16943 15265 16946
rect 15420 16946 15426 18482
rect 15460 16946 15466 18482
rect 15508 18482 15554 18494
rect 15508 17857 15514 18482
rect 15506 17601 15514 17857
rect 15098 16934 15144 16943
rect 15420 16934 15466 16946
rect 15508 16946 15514 17601
rect 15548 17857 15554 18482
rect 16253 18409 16270 18537
rect 15787 17870 15974 18232
rect 16264 18140 16270 18409
rect 16308 18409 16326 18537
rect 16308 18140 16314 18409
rect 16788 18350 16878 18352
rect 16264 18128 16314 18140
rect 16780 18346 16880 18350
rect 16780 18280 16800 18346
rect 16866 18280 16880 18346
rect 16780 18040 16880 18280
rect 16780 17940 16790 18040
rect 16870 17940 16880 18040
rect 16780 17930 16880 17940
rect 17330 18040 17530 18060
rect 15780 17857 16980 17870
rect 15548 17836 16980 17857
rect 15548 17601 15878 17836
rect 15548 16946 15554 17601
rect 15872 17439 15878 17601
rect 15916 17610 16980 17836
rect 17330 17740 17350 18040
rect 17510 17740 17530 18040
rect 17330 17720 17412 17740
rect 15916 17602 15974 17610
rect 15916 17601 15934 17602
rect 15916 17439 15922 17601
rect 15872 17427 15922 17439
rect 16720 17530 16980 17610
rect 15872 17305 15922 17317
rect 15872 16984 15878 17305
rect 15508 16934 15554 16946
rect 14596 16434 14756 16908
rect 15816 16908 15878 16984
rect 15916 16984 15922 17305
rect 16264 17306 16314 17318
rect 16264 17141 16270 17306
rect 15916 16908 15976 16984
rect 14596 16334 14616 16434
rect 14736 16334 14756 16434
rect 14596 16314 14756 16334
rect 15016 16899 15126 16904
rect 15016 16896 15130 16899
rect 15016 16862 15060 16896
rect 15094 16862 15130 16896
rect 15016 16484 15130 16862
rect 15444 16896 15533 16905
rect 15444 16862 15470 16896
rect 15504 16862 15533 16896
rect 15444 16692 15533 16862
rect 15444 16566 15456 16692
rect 15515 16566 15533 16692
rect 15444 16554 15533 16566
rect 13516 16279 14484 16289
rect 15016 16284 15026 16484
rect 15116 16284 15130 16484
rect 15816 16434 15976 16908
rect 16249 16909 16270 17141
rect 16308 17141 16314 17306
rect 16720 17300 16760 17530
rect 16950 17300 16980 17530
rect 17406 17524 17412 17720
rect 17450 17720 17530 17740
rect 17450 17524 17456 17720
rect 17406 17512 17456 17524
rect 16720 17270 16980 17300
rect 16308 16909 18052 17141
rect 16249 16884 18052 16909
rect 15816 16334 15836 16434
rect 15946 16334 15976 16434
rect 15816 16308 15976 16334
rect 15016 16274 15130 16284
rect 13000 16104 16242 16224
rect 13572 15536 13692 16104
rect 14742 16004 14842 16014
rect 14742 15984 14752 16004
rect 14552 15976 14752 15984
rect 14832 15984 14842 16004
rect 14832 15976 15192 15984
rect 14552 15942 14566 15976
rect 14600 15944 14752 15976
rect 14832 15944 14950 15976
rect 14600 15942 14758 15944
rect 14792 15942 14950 15944
rect 14984 15942 15142 15976
rect 15176 15942 15192 15976
rect 14552 15934 15192 15942
rect 16122 15946 16242 16104
rect 17212 16024 17292 16044
rect 17212 15990 17236 16024
rect 17270 15990 17292 16024
rect 17212 15984 17292 15990
rect 13572 15502 13616 15536
rect 13650 15502 13692 15536
rect 13572 15494 13692 15502
rect 14416 15892 14462 15904
rect 13566 15452 13612 15464
rect 13507 15439 13572 15452
rect 13507 15320 13520 15439
rect 13507 15307 13572 15320
rect 13566 14020 13572 15307
rect 13480 13916 13572 14020
rect 13606 13916 13612 15452
rect 13480 13904 13612 13916
rect 13654 15452 13700 15464
rect 13654 13916 13660 15452
rect 13694 13916 13700 15452
rect 14416 14034 14422 15892
rect 13654 13904 13700 13916
rect 14413 13916 14422 14034
rect 14456 14034 14462 15892
rect 14493 15894 14563 15904
rect 14493 15794 14502 15894
rect 14554 15794 14563 15894
rect 14493 15784 14518 15794
rect 14456 14024 14483 14034
rect 14474 13924 14483 14024
rect 14456 13916 14483 13924
rect 14413 13914 14483 13916
rect 14512 13916 14518 15784
rect 14552 15784 14563 15794
rect 14608 15892 14654 15904
rect 14552 13916 14558 15784
rect 14608 14034 14614 15892
rect 14416 13904 14462 13914
rect 14512 13904 14558 13916
rect 14593 14024 14614 14034
rect 14648 14034 14654 15892
rect 14693 15894 14763 15904
rect 14693 15794 14702 15894
rect 14754 15794 14763 15894
rect 14693 15784 14710 15794
rect 14648 14024 14663 14034
rect 14593 13924 14602 14024
rect 14654 13924 14663 14024
rect 14593 13916 14614 13924
rect 14648 13916 14663 13924
rect 14593 13914 14663 13916
rect 14704 13916 14710 15784
rect 14744 15784 14763 15794
rect 14800 15892 14846 15904
rect 14744 13916 14750 15784
rect 14800 14034 14806 15892
rect 14608 13904 14654 13914
rect 14704 13904 14750 13916
rect 14783 14024 14806 14034
rect 14840 14034 14846 15892
rect 14883 15894 14953 15904
rect 14883 15794 14892 15894
rect 14944 15794 14953 15894
rect 14883 15784 14902 15794
rect 14840 14024 14853 14034
rect 14783 13924 14792 14024
rect 14844 13924 14853 14024
rect 14783 13916 14806 13924
rect 14840 13916 14853 13924
rect 14783 13914 14853 13916
rect 14896 13916 14902 15784
rect 14936 15784 14953 15794
rect 14992 15892 15038 15904
rect 14936 13916 14942 15784
rect 14992 14034 14998 15892
rect 14800 13904 14846 13914
rect 14896 13904 14942 13916
rect 14973 14024 14998 14034
rect 15032 14034 15038 15892
rect 15073 15894 15143 15904
rect 15073 15794 15082 15894
rect 15134 15794 15143 15894
rect 15073 15784 15094 15794
rect 15032 14024 15043 14034
rect 14973 13924 14982 14024
rect 15034 13924 15043 14024
rect 14973 13916 14998 13924
rect 15032 13916 15043 13924
rect 14973 13914 15043 13916
rect 15088 13916 15094 15784
rect 15128 15784 15143 15794
rect 15184 15892 15230 15904
rect 15128 13916 15134 15784
rect 15184 14034 15190 15892
rect 14992 13904 15038 13914
rect 15088 13904 15134 13916
rect 15163 14024 15190 14034
rect 15224 14034 15230 15892
rect 16122 15549 16164 15946
rect 16202 15549 16242 15946
rect 16122 15524 16242 15549
rect 17086 15931 17132 15943
rect 16122 14275 16242 14314
rect 15163 13924 15172 14024
rect 15163 13916 15190 13924
rect 15224 13916 15233 14034
rect 15163 13914 15233 13916
rect 15184 13904 15230 13914
rect 13480 13195 13572 13904
rect 16122 13878 16164 14275
rect 16202 13878 16242 14275
rect 17086 14064 17092 15931
rect 17073 14054 17092 14064
rect 17126 14064 17132 15931
rect 17173 15934 17243 15944
rect 17173 15834 17182 15934
rect 17234 15834 17243 15934
rect 17173 15824 17188 15834
rect 17126 14054 17143 14064
rect 17073 13954 17082 14054
rect 17134 13954 17143 14054
rect 17073 13944 17143 13954
rect 17182 13955 17188 15824
rect 17222 15824 17243 15834
rect 17278 15931 17324 15943
rect 17222 13955 17228 15824
rect 17278 14064 17284 15931
rect 17086 13943 17132 13944
rect 17182 13943 17228 13955
rect 17273 14054 17284 14064
rect 17318 14064 17324 15931
rect 17363 15934 17433 15944
rect 17363 15834 17372 15934
rect 17424 15834 17433 15934
rect 17363 15824 17380 15834
rect 17318 14054 17343 14064
rect 17273 13954 17282 14054
rect 17334 13954 17343 14054
rect 17273 13944 17343 13954
rect 17374 13955 17380 15824
rect 17414 15824 17433 15834
rect 17414 13955 17420 15824
rect 17278 13943 17324 13944
rect 17374 13943 17420 13955
rect 17122 13913 17382 13914
rect 13604 13871 13662 13872
rect 13600 13866 13668 13871
rect 13600 13864 13616 13866
rect 13650 13864 13668 13866
rect 13600 13813 13611 13864
rect 13601 13803 13611 13813
rect 13663 13803 13668 13864
rect 14452 13866 15092 13874
rect 14452 13832 14470 13866
rect 14504 13832 14662 13866
rect 14696 13832 14854 13866
rect 14888 13832 15046 13866
rect 15080 13832 15092 13866
rect 14452 13824 15092 13832
rect 13601 13794 13668 13803
rect 16122 13354 16242 13878
rect 17000 13896 17385 13913
rect 17000 13862 17140 13896
rect 17174 13862 17332 13896
rect 17366 13862 17385 13896
rect 17000 13795 17385 13862
rect 16112 13344 16252 13354
rect 16112 13284 16132 13344
rect 16232 13284 16252 13344
rect 16112 13264 16252 13284
rect 17000 13313 17118 13795
rect 17000 13273 17021 13313
rect 17093 13273 17118 13313
rect 17000 13254 17118 13273
rect 13480 13133 13500 13195
rect 13552 13133 13572 13195
rect 13480 13116 13572 13133
rect 13603 13173 13824 13219
rect 13480 13115 13571 13116
rect 13603 13070 13649 13173
rect 13778 13070 13824 13173
rect 13959 13170 14180 13216
rect 13959 13070 14005 13170
rect 14134 13070 14180 13170
rect 14312 13175 14533 13221
rect 14312 13070 14358 13175
rect 14487 13070 14533 13175
rect 14660 13167 14881 13213
rect 13428 13058 13474 13070
rect 13516 13062 13562 13070
rect 13428 11082 13434 13058
rect 13468 11082 13474 13058
rect 13508 13058 13570 13062
rect 13508 13052 13522 13058
rect 13556 13052 13570 13058
rect 13508 12960 13512 13052
rect 13566 12960 13570 13052
rect 13603 13058 13650 13070
rect 13692 13068 13738 13070
rect 13603 13051 13610 13058
rect 13508 12950 13522 12960
rect 13428 10970 13474 11082
rect 13516 11082 13522 12950
rect 13556 12950 13570 12960
rect 13556 11082 13562 12950
rect 13604 11101 13610 13051
rect 13516 11070 13562 11082
rect 13603 11082 13610 11101
rect 13644 11082 13650 13058
rect 13678 13058 13743 13068
rect 13678 13055 13698 13058
rect 13732 13055 13743 13058
rect 13678 12966 13685 13055
rect 13737 12966 13743 13055
rect 13778 13058 13826 13070
rect 13868 13062 13914 13070
rect 13778 13042 13786 13058
rect 13678 12954 13698 12966
rect 13603 11070 13650 11082
rect 13692 11082 13698 12954
rect 13732 12954 13743 12966
rect 13732 11082 13738 12954
rect 13692 11070 13738 11082
rect 13780 11082 13786 13042
rect 13820 11090 13826 13058
rect 13856 13058 13918 13062
rect 13856 13052 13874 13058
rect 13908 13052 13918 13058
rect 13856 12960 13860 13052
rect 13914 12960 13918 13052
rect 13856 12950 13874 12960
rect 13820 11082 13827 11090
rect 13780 11070 13827 11082
rect 13868 11082 13874 12950
rect 13908 12950 13918 12960
rect 13956 13058 14005 13070
rect 13908 11082 13914 12950
rect 13868 11070 13914 11082
rect 13956 11082 13962 13058
rect 13996 13048 14005 13058
rect 14035 13058 14100 13070
rect 14035 13057 14050 13058
rect 14084 13057 14100 13058
rect 13996 11082 14002 13048
rect 14035 12968 14042 13057
rect 14094 12968 14100 13057
rect 14035 12956 14050 12968
rect 13603 10970 13649 11070
rect 13428 10924 13649 10970
rect 13781 10968 13827 11070
rect 13956 10968 14002 11082
rect 14044 11082 14050 12956
rect 14084 12956 14100 12968
rect 14132 13058 14180 13070
rect 14220 13068 14266 13070
rect 14084 11082 14090 12956
rect 14044 11070 14090 11082
rect 14132 11082 14138 13058
rect 14172 13039 14180 13058
rect 14212 13058 14274 13068
rect 14172 11082 14178 13039
rect 14212 12966 14216 13058
rect 14270 12966 14274 13058
rect 14212 12956 14226 12966
rect 13781 10922 14002 10968
rect 14132 10970 14178 11082
rect 14220 11082 14226 12956
rect 14260 12956 14274 12966
rect 14308 13058 14358 13070
rect 14260 11082 14266 12956
rect 14308 11101 14314 13058
rect 14220 11070 14266 11082
rect 14307 11082 14314 11101
rect 14348 13053 14358 13058
rect 14388 13058 14453 13070
rect 14388 13057 14402 13058
rect 14436 13057 14453 13058
rect 14348 11082 14354 13053
rect 14388 12968 14395 13057
rect 14447 12968 14453 13057
rect 14388 12956 14402 12968
rect 14307 11070 14354 11082
rect 14396 11082 14402 12956
rect 14436 12956 14453 12968
rect 14484 13058 14533 13070
rect 14572 13066 14618 13070
rect 14436 11082 14442 12956
rect 14396 11070 14442 11082
rect 14484 11082 14490 13058
rect 14524 13044 14533 13058
rect 14562 13058 14624 13066
rect 14562 13056 14578 13058
rect 14612 13056 14624 13058
rect 14524 11082 14530 13044
rect 14562 12964 14566 13056
rect 14620 12964 14624 13056
rect 14562 12954 14578 12964
rect 14307 10970 14353 11070
rect 14484 10994 14530 11082
rect 14572 11082 14578 12954
rect 14612 12954 14624 12964
rect 14660 13058 14706 13167
rect 14612 11082 14618 12954
rect 14660 11101 14666 13058
rect 14572 11070 14618 11082
rect 14659 11082 14666 11101
rect 14700 11082 14706 13058
rect 14740 13058 14805 13071
rect 14740 12969 14747 13058
rect 14799 12969 14805 13058
rect 14835 13070 14881 13167
rect 15016 13175 15237 13221
rect 15016 13070 15062 13175
rect 15191 13070 15237 13175
rect 15366 13175 15587 13221
rect 15366 13070 15412 13175
rect 15541 13070 15587 13175
rect 15720 13173 15941 13219
rect 15720 13070 15766 13173
rect 15895 13070 15941 13173
rect 16069 13171 16290 13217
rect 16069 13070 16115 13171
rect 14835 13058 14882 13070
rect 14924 13066 14970 13070
rect 14835 13036 14842 13058
rect 14740 12957 14754 12969
rect 14659 11070 14706 11082
rect 14748 11082 14754 12957
rect 14788 12957 14805 12969
rect 14788 11082 14794 12957
rect 14748 11070 14794 11082
rect 14836 11082 14842 13036
rect 14876 11092 14882 13058
rect 14916 13058 14978 13066
rect 14916 13056 14930 13058
rect 14964 13056 14978 13058
rect 14916 12964 14920 13056
rect 14974 12964 14978 13056
rect 14916 12954 14930 12964
rect 14876 11082 14883 11092
rect 14836 11070 14883 11082
rect 14924 11082 14930 12954
rect 14964 12954 14978 12964
rect 15012 13058 15062 13070
rect 14964 11082 14970 12954
rect 14924 11070 14970 11082
rect 15012 11082 15018 13058
rect 15052 13053 15062 13058
rect 15091 13058 15156 13070
rect 15091 13057 15106 13058
rect 15140 13057 15156 13058
rect 15052 11082 15058 13053
rect 15091 12968 15098 13057
rect 15150 12968 15156 13057
rect 15091 12956 15106 12968
rect 14659 10994 14705 11070
rect 14132 10924 14353 10970
rect 14482 10924 14705 10994
rect 14837 10970 14883 11070
rect 15012 10970 15058 11082
rect 15100 11082 15106 12956
rect 15140 12956 15156 12968
rect 15188 13058 15237 13070
rect 15276 13068 15322 13070
rect 15140 11082 15146 12956
rect 15100 11070 15146 11082
rect 15188 11082 15194 13058
rect 15228 13044 15237 13058
rect 15270 13058 15332 13068
rect 15228 11092 15234 13044
rect 15270 12966 15274 13058
rect 15328 12966 15332 13058
rect 15270 12956 15282 12966
rect 15228 11082 15236 11092
rect 15188 11070 15236 11082
rect 15276 11082 15282 12956
rect 15316 12956 15332 12966
rect 15364 13058 15412 13070
rect 15452 13065 15498 13070
rect 15316 11082 15322 12956
rect 15276 11070 15322 11082
rect 15364 11082 15370 13058
rect 15404 13053 15412 13058
rect 15443 13058 15508 13065
rect 15404 11101 15410 13053
rect 15443 13052 15458 13058
rect 15492 13052 15508 13058
rect 15443 12963 15450 13052
rect 15502 12963 15508 13052
rect 15443 12951 15458 12963
rect 15404 11082 15411 11101
rect 15364 11070 15411 11082
rect 15452 11082 15458 12951
rect 15492 12951 15508 12963
rect 15540 13058 15587 13070
rect 15628 13068 15674 13070
rect 15492 11082 15498 12951
rect 15452 11070 15498 11082
rect 15540 11082 15546 13058
rect 15580 13044 15587 13058
rect 15622 13058 15684 13068
rect 15580 11082 15586 13044
rect 15622 12966 15626 13058
rect 15680 12966 15684 13058
rect 15622 12956 15634 12966
rect 14837 10924 15058 10970
rect 15190 10970 15236 11070
rect 15365 10970 15411 11070
rect 15190 10924 15411 10970
rect 15540 10971 15586 11082
rect 15628 11082 15634 12956
rect 15668 12956 15684 12966
rect 15716 13058 15766 13070
rect 15804 13065 15850 13070
rect 15668 11082 15674 12956
rect 15716 11102 15722 13058
rect 15628 11070 15674 11082
rect 15715 11082 15722 11102
rect 15756 13051 15766 13058
rect 15796 13058 15861 13065
rect 15796 13052 15810 13058
rect 15844 13052 15861 13058
rect 15756 11082 15762 13051
rect 15796 12963 15803 13052
rect 15855 12963 15861 13052
rect 15796 12951 15810 12963
rect 15715 11070 15762 11082
rect 15804 11082 15810 12951
rect 15844 12951 15861 12963
rect 15892 13058 15941 13070
rect 15980 13064 16026 13070
rect 15844 11082 15850 12951
rect 15804 11070 15850 11082
rect 15892 11082 15898 13058
rect 15932 13042 15941 13058
rect 15972 13058 16034 13064
rect 15972 13054 15986 13058
rect 16020 13054 16034 13058
rect 15932 11093 15938 13042
rect 15972 12962 15976 13054
rect 16030 12962 16034 13054
rect 15972 12952 15986 12962
rect 15932 11082 15941 11093
rect 15892 11070 15941 11082
rect 15980 11082 15986 12952
rect 16020 12952 16034 12962
rect 16068 13058 16115 13070
rect 16156 13065 16202 13070
rect 16020 11082 16026 12952
rect 15980 11070 16026 11082
rect 16068 11082 16074 13058
rect 16108 13049 16115 13058
rect 16148 13058 16213 13065
rect 16148 13052 16162 13058
rect 16196 13052 16213 13058
rect 16108 11102 16114 13049
rect 16148 12963 16155 13052
rect 16207 12963 16213 13052
rect 16148 12951 16162 12963
rect 16108 11082 16116 11102
rect 16068 11070 16116 11082
rect 16156 11082 16162 12951
rect 16196 12951 16213 12963
rect 16244 13058 16290 13171
rect 16423 13175 16644 13221
rect 16423 13070 16469 13175
rect 16598 13070 16644 13175
rect 16777 13171 16998 13217
rect 16777 13070 16823 13171
rect 16952 13070 16998 13171
rect 17130 13171 17351 13217
rect 17130 13070 17176 13171
rect 17305 13070 17351 13171
rect 16332 13064 16378 13070
rect 16196 11082 16202 12951
rect 16156 11070 16202 11082
rect 16244 11082 16250 13058
rect 16284 11082 16290 13058
rect 16326 13058 16388 13064
rect 16326 13054 16338 13058
rect 16372 13054 16388 13058
rect 16326 12962 16330 13054
rect 16384 12962 16388 13054
rect 16326 12952 16338 12962
rect 15715 10971 15761 11070
rect 15540 10925 15761 10971
rect 15895 10971 15941 11070
rect 16070 10971 16116 11070
rect 15895 10925 16116 10971
rect 16244 10971 16290 11082
rect 16332 11082 16338 12952
rect 16372 12952 16388 12962
rect 16420 13058 16469 13070
rect 16508 13064 16554 13070
rect 16372 11082 16378 12952
rect 16420 11102 16426 13058
rect 16332 11070 16378 11082
rect 16419 11082 16426 11102
rect 16460 13053 16469 13058
rect 16502 13058 16567 13064
rect 16460 11082 16466 13053
rect 16502 13051 16514 13058
rect 16548 13051 16567 13058
rect 16502 12962 16509 13051
rect 16561 12962 16567 13051
rect 16502 12950 16514 12962
rect 16419 11070 16466 11082
rect 16508 11082 16514 12950
rect 16548 12950 16567 12962
rect 16596 13058 16644 13070
rect 16684 13066 16730 13070
rect 16548 11082 16554 12950
rect 16508 11070 16554 11082
rect 16596 11082 16602 13058
rect 16636 13044 16644 13058
rect 16676 13058 16738 13066
rect 16676 13056 16690 13058
rect 16724 13056 16738 13058
rect 16636 11082 16642 13044
rect 16676 12964 16680 13056
rect 16734 12964 16738 13056
rect 16676 12954 16690 12964
rect 16419 10971 16465 11070
rect 16244 10925 16465 10971
rect 16596 10970 16642 11082
rect 16684 11082 16690 12954
rect 16724 12954 16738 12964
rect 16772 13058 16823 13070
rect 16724 11082 16730 12954
rect 16772 11101 16778 13058
rect 16684 11070 16730 11082
rect 16771 11082 16778 11101
rect 16812 13049 16823 13058
rect 16851 13058 16916 13070
rect 16851 13057 16866 13058
rect 16900 13057 16916 13058
rect 16812 11082 16818 13049
rect 16851 12968 16858 13057
rect 16910 12968 16916 13057
rect 16851 12956 16866 12968
rect 16771 11070 16818 11082
rect 16860 11082 16866 12956
rect 16900 12956 16916 12968
rect 16948 13058 16998 13070
rect 17036 13066 17082 13070
rect 16900 11082 16906 12956
rect 16860 11070 16906 11082
rect 16948 11082 16954 13058
rect 16988 13040 16998 13058
rect 17030 13058 17092 13066
rect 17030 13056 17042 13058
rect 17076 13056 17092 13058
rect 16988 11082 16994 13040
rect 17030 12964 17034 13056
rect 17088 12964 17092 13056
rect 17030 12954 17042 12964
rect 16771 10970 16817 11070
rect 16596 10924 16817 10970
rect 16948 10971 16994 11082
rect 17036 11082 17042 12954
rect 17076 12954 17092 12964
rect 17124 13058 17176 13070
rect 17212 13065 17258 13070
rect 17076 11082 17082 12954
rect 17124 11102 17130 13058
rect 17036 11070 17082 11082
rect 17123 11082 17130 11102
rect 17164 13049 17176 13058
rect 17204 13058 17269 13065
rect 17204 13052 17218 13058
rect 17252 13052 17269 13058
rect 17164 11082 17170 13049
rect 17204 12963 17211 13052
rect 17263 12963 17269 13052
rect 17204 12951 17218 12963
rect 17123 11070 17170 11082
rect 17212 11082 17218 12951
rect 17252 12951 17269 12963
rect 17300 13058 17351 13070
rect 17252 11082 17258 12951
rect 17212 11070 17258 11082
rect 17300 11082 17306 13058
rect 17340 13040 17351 13058
rect 17381 13058 17446 13070
rect 17381 13057 17394 13058
rect 17428 13057 17446 13058
rect 17340 11093 17346 13040
rect 17381 12968 17388 13057
rect 17440 12968 17446 13057
rect 17381 12956 17394 12968
rect 17340 11082 17347 11093
rect 17300 11070 17347 11082
rect 17388 11082 17394 12956
rect 17428 12956 17446 12968
rect 17476 13058 17522 13070
rect 17428 11082 17434 12956
rect 17388 11070 17434 11082
rect 17476 11082 17482 13058
rect 17516 11082 17522 13058
rect 17123 10971 17169 11070
rect 16948 10925 17169 10971
rect 17301 10971 17347 11070
rect 17476 10971 17522 11082
rect 17301 10925 17522 10971
rect 13467 10874 13597 10886
rect 13467 10815 13482 10874
rect 13581 10815 13597 10874
rect 13467 10368 13597 10815
rect 14482 10714 14702 10924
rect 17342 10874 17482 10894
rect 17342 10784 17362 10874
rect 17462 10784 17482 10874
rect 14482 10654 14502 10714
rect 14682 10654 14702 10714
rect 14482 10634 14702 10654
rect 17264 10624 17570 10784
rect 17264 10372 17276 10624
rect 17542 10372 17570 10624
rect 17264 10356 17570 10372
rect 17795 10640 18052 16884
rect 17795 10380 17806 10640
rect 18034 10380 18052 10640
rect 17795 10364 18052 10380
rect 4162 9718 26614 9766
rect 4162 8388 4218 9718
rect 5576 9698 26614 9718
rect 5576 9688 25266 9698
rect 5576 8938 13906 9688
rect 16938 8938 25266 9688
rect 5576 8388 25266 8938
rect 4162 8378 25266 8388
rect 26538 8378 26614 9698
rect 4162 8342 26614 8378
rect 2149 7480 28685 7576
rect 2149 6346 2324 7480
rect 3678 7470 28685 7480
rect 3678 6346 27174 7470
rect 2149 6336 27174 6346
rect 28528 6336 28685 7470
rect 2149 6246 28685 6336
<< via1 >>
rect 2340 27686 3694 28820
rect 27180 27758 28534 28892
rect 4246 25634 5518 26954
rect 25304 25642 26576 26962
rect 16820 24600 16900 24610
rect 16820 24562 16892 24600
rect 16892 24562 16900 24600
rect 16820 24520 16900 24562
rect 13664 23042 13792 23372
rect 15272 23364 15414 23612
rect 16290 23430 16430 23560
rect 12559 17700 12791 17968
rect 14050 23050 14066 23132
rect 14066 23050 14100 23132
rect 14100 23050 14102 23132
rect 13960 21170 13970 21252
rect 13970 21170 14004 21252
rect 14004 21170 14012 21252
rect 14250 23050 14258 23132
rect 14258 23050 14292 23132
rect 14292 23050 14302 23132
rect 14150 21170 14162 21252
rect 14162 21170 14196 21252
rect 14196 21170 14202 21252
rect 14440 23050 14450 23132
rect 14450 23050 14484 23132
rect 14484 23050 14492 23132
rect 14340 21170 14354 21252
rect 14354 21170 14388 21252
rect 14388 21170 14392 21252
rect 14630 23050 14642 23132
rect 14642 23050 14676 23132
rect 14676 23050 14682 23132
rect 14530 21170 14546 21252
rect 14546 21170 14580 21252
rect 14580 21170 14582 21252
rect 14830 23040 14900 23140
rect 14730 21170 14738 21252
rect 14738 21170 14772 21252
rect 14772 21170 14782 21252
rect 15910 23090 15926 23172
rect 15926 23090 15960 23172
rect 15960 23090 15962 23172
rect 15810 21210 15830 21292
rect 15830 21210 15862 21292
rect 16100 23090 16118 23172
rect 16118 23090 16152 23172
rect 16010 21210 16022 21292
rect 16022 21210 16056 21292
rect 16056 21210 16062 21292
rect 16750 24028 16803 24031
rect 16750 23920 16758 24028
rect 16758 23920 16792 24028
rect 16792 23920 16803 24028
rect 16658 22052 16662 22160
rect 16662 22052 16696 22160
rect 16696 22052 16711 22160
rect 16658 22049 16711 22052
rect 16940 24028 16993 24031
rect 16940 23920 16950 24028
rect 16950 23920 16984 24028
rect 16984 23920 16993 24028
rect 16839 22052 16854 22160
rect 16854 22052 16888 22160
rect 16888 22052 16892 22160
rect 16839 22049 16892 22052
rect 17130 24028 17183 24031
rect 17130 23920 17142 24028
rect 17142 23920 17176 24028
rect 17176 23920 17183 24028
rect 17029 22052 17046 22160
rect 17046 22052 17080 22160
rect 17080 22052 17082 22160
rect 17029 22049 17082 22052
rect 17320 24028 17373 24031
rect 17320 23920 17334 24028
rect 17334 23920 17368 24028
rect 17368 23920 17373 24028
rect 17220 22052 17238 22163
rect 17238 22052 17272 22163
rect 17272 22052 17273 22163
rect 17520 24028 17573 24031
rect 17520 23920 17526 24028
rect 17526 23920 17560 24028
rect 17560 23920 17573 24028
rect 17419 22052 17430 22161
rect 17430 22052 17464 22161
rect 17464 22052 17472 22161
rect 17419 22050 17472 22052
rect 17610 22052 17622 22162
rect 17622 22052 17656 22162
rect 17656 22052 17663 22162
rect 17610 22051 17663 22052
rect 16864 20932 17006 21322
rect 14920 20518 15460 20550
rect 14920 20490 14974 20518
rect 14974 20490 15008 20518
rect 15008 20490 15166 20518
rect 15166 20490 15200 20518
rect 15200 20490 15358 20518
rect 15358 20490 15392 20518
rect 15392 20490 15460 20518
rect 14910 20320 14926 20430
rect 14926 20320 14960 20430
rect 14960 20320 14970 20430
rect 14820 19180 14830 19290
rect 14830 19180 14864 19290
rect 14864 19180 14880 19290
rect 15100 20320 15118 20430
rect 15118 20320 15152 20430
rect 15152 20320 15160 20430
rect 15010 19180 15022 19290
rect 15022 19180 15056 19290
rect 15056 19180 15070 19290
rect 15300 20320 15310 20430
rect 15310 20320 15344 20430
rect 15344 20320 15360 20430
rect 15200 19180 15214 19290
rect 15214 19180 15248 19290
rect 15248 19180 15260 19290
rect 15490 20320 15502 20430
rect 15502 20320 15536 20430
rect 15536 20320 15550 20430
rect 15390 19180 15406 19290
rect 15406 19180 15440 19290
rect 15440 19180 15450 19290
rect 16070 19948 16130 19950
rect 16070 19840 16086 19948
rect 16086 19840 16120 19948
rect 16120 19840 16130 19948
rect 15970 19172 15990 19280
rect 15990 19172 16024 19280
rect 16024 19172 16030 19280
rect 15970 19170 16030 19172
rect 16260 19948 16320 19950
rect 16260 19840 16278 19948
rect 16278 19840 16312 19948
rect 16312 19840 16320 19948
rect 16170 19172 16182 19280
rect 16182 19172 16216 19280
rect 16216 19172 16230 19280
rect 16170 19170 16230 19172
rect 16500 19030 16600 19120
rect 17040 19170 17210 19260
rect 14156 16574 14286 16694
rect 14654 17606 14658 17833
rect 14658 17606 14696 17833
rect 14696 17606 14737 17833
rect 13528 16289 13592 16384
rect 15115 17606 15138 17835
rect 15138 17606 15175 17835
rect 16790 17940 16870 18040
rect 17350 17921 17510 18040
rect 17350 17740 17412 17921
rect 17412 17740 17450 17921
rect 17450 17740 17510 17921
rect 15456 16566 15515 16692
rect 15026 16284 15116 16484
rect 16760 17300 16950 17530
rect 14752 15976 14832 16004
rect 14752 15944 14758 15976
rect 14758 15944 14792 15976
rect 14792 15944 14832 15976
rect 13520 15320 13572 15439
rect 13572 15320 13589 15439
rect 14502 15892 14554 15894
rect 14502 15794 14518 15892
rect 14518 15794 14552 15892
rect 14552 15794 14554 15892
rect 14422 13924 14456 14024
rect 14456 13924 14474 14024
rect 14702 15892 14754 15894
rect 14702 15794 14710 15892
rect 14710 15794 14744 15892
rect 14744 15794 14754 15892
rect 14602 13924 14614 14024
rect 14614 13924 14648 14024
rect 14648 13924 14654 14024
rect 14892 15892 14944 15894
rect 14892 15794 14902 15892
rect 14902 15794 14936 15892
rect 14936 15794 14944 15892
rect 14792 13924 14806 14024
rect 14806 13924 14840 14024
rect 14840 13924 14844 14024
rect 15082 15892 15134 15894
rect 15082 15794 15094 15892
rect 15094 15794 15128 15892
rect 15128 15794 15134 15892
rect 14982 13924 14998 14024
rect 14998 13924 15032 14024
rect 15032 13924 15034 14024
rect 15172 13924 15190 14024
rect 15190 13924 15224 14024
rect 17182 15931 17234 15934
rect 17182 15834 17188 15931
rect 17188 15834 17222 15931
rect 17222 15834 17234 15931
rect 17082 13955 17092 14054
rect 17092 13955 17126 14054
rect 17126 13955 17134 14054
rect 17082 13954 17134 13955
rect 17372 15931 17424 15934
rect 17372 15834 17380 15931
rect 17380 15834 17414 15931
rect 17414 15834 17424 15931
rect 17282 13955 17284 14054
rect 17284 13955 17318 14054
rect 17318 13955 17334 14054
rect 17282 13954 17334 13955
rect 13611 13832 13616 13864
rect 13616 13832 13650 13864
rect 13650 13832 13663 13864
rect 13611 13803 13663 13832
rect 13512 12960 13522 13052
rect 13522 12960 13556 13052
rect 13556 12960 13566 13052
rect 13685 12966 13698 13055
rect 13698 12966 13732 13055
rect 13732 12966 13737 13055
rect 13860 12960 13874 13052
rect 13874 12960 13908 13052
rect 13908 12960 13914 13052
rect 14042 12968 14050 13057
rect 14050 12968 14084 13057
rect 14084 12968 14094 13057
rect 14216 12966 14226 13058
rect 14226 12966 14260 13058
rect 14260 12966 14270 13058
rect 14395 12968 14402 13057
rect 14402 12968 14436 13057
rect 14436 12968 14447 13057
rect 14566 12964 14578 13056
rect 14578 12964 14612 13056
rect 14612 12964 14620 13056
rect 14747 12969 14754 13058
rect 14754 12969 14788 13058
rect 14788 12969 14799 13058
rect 14920 12964 14930 13056
rect 14930 12964 14964 13056
rect 14964 12964 14974 13056
rect 15098 12968 15106 13057
rect 15106 12968 15140 13057
rect 15140 12968 15150 13057
rect 15274 12966 15282 13058
rect 15282 12966 15316 13058
rect 15316 12966 15328 13058
rect 15450 12963 15458 13052
rect 15458 12963 15492 13052
rect 15492 12963 15502 13052
rect 15626 12966 15634 13058
rect 15634 12966 15668 13058
rect 15668 12966 15680 13058
rect 15803 12963 15810 13052
rect 15810 12963 15844 13052
rect 15844 12963 15855 13052
rect 15976 12962 15986 13054
rect 15986 12962 16020 13054
rect 16020 12962 16030 13054
rect 16155 12963 16162 13052
rect 16162 12963 16196 13052
rect 16196 12963 16207 13052
rect 16330 12962 16338 13054
rect 16338 12962 16372 13054
rect 16372 12962 16384 13054
rect 16509 12962 16514 13051
rect 16514 12962 16548 13051
rect 16548 12962 16561 13051
rect 16680 12964 16690 13056
rect 16690 12964 16724 13056
rect 16724 12964 16734 13056
rect 16858 12968 16866 13057
rect 16866 12968 16900 13057
rect 16900 12968 16910 13057
rect 17034 12964 17042 13056
rect 17042 12964 17076 13056
rect 17076 12964 17088 13056
rect 17211 12963 17218 13052
rect 17218 12963 17252 13052
rect 17252 12963 17263 13052
rect 17388 12968 17394 13057
rect 17394 12968 17428 13057
rect 17428 12968 17440 13057
rect 17276 10372 17542 10624
rect 17806 10380 18034 10640
rect 4218 8388 5576 9718
rect 25266 8378 26538 9698
rect 2324 6346 3678 7480
rect 27174 6336 28528 7470
<< metal2 >>
rect 2168 28820 3820 28952
rect 2168 27686 2340 28820
rect 3694 27686 3820 28820
rect 2168 7480 3820 27686
rect 27052 28892 28704 28952
rect 27052 27758 27180 28892
rect 28534 27758 28704 28892
rect 4162 26954 5612 26992
rect 4162 25634 4246 26954
rect 5518 25634 5612 26954
rect 4162 9718 5612 25634
rect 25230 26962 26614 27010
rect 25230 25642 25304 26962
rect 26576 25642 26614 26962
rect 17828 25332 18030 25342
rect 12324 25304 12582 25328
rect 12324 24874 12340 25304
rect 12564 24874 12582 25304
rect 12324 23390 12582 24874
rect 17828 25110 17844 25332
rect 18020 25110 18030 25332
rect 16810 24610 16910 24620
rect 16810 24520 16820 24610
rect 16900 24520 16910 24610
rect 16810 24426 16910 24520
rect 17828 24426 18030 25110
rect 16810 24250 18030 24426
rect 16810 24050 16910 24250
rect 17828 24248 18030 24250
rect 18170 25302 18480 25326
rect 18170 25024 18192 25302
rect 18456 25024 18480 25302
rect 16810 24041 16950 24050
rect 16743 24040 17003 24041
rect 17123 24040 17193 24041
rect 17313 24040 17383 24041
rect 17513 24040 17583 24041
rect 16740 24031 17583 24040
rect 16740 23920 16750 24031
rect 16803 23920 16940 24031
rect 16993 23920 17130 24031
rect 17183 23920 17320 24031
rect 17373 23920 17520 24031
rect 17573 23920 17583 24031
rect 16740 23911 17583 23920
rect 16740 23910 17570 23911
rect 15260 23612 15432 23632
rect 12324 23388 13786 23390
rect 12324 23372 13802 23388
rect 12324 23042 13664 23372
rect 13792 23042 13802 23372
rect 15260 23364 15272 23612
rect 15414 23364 15432 23612
rect 16270 23560 16450 23580
rect 16270 23430 16290 23560
rect 16430 23430 16450 23560
rect 16270 23410 16450 23430
rect 15260 23312 15432 23364
rect 15901 23190 15971 23191
rect 16091 23190 16161 23191
rect 15901 23172 16161 23190
rect 12324 23032 13802 23042
rect 12334 23030 13802 23032
rect 14041 23150 14111 23151
rect 14241 23150 14311 23151
rect 14431 23150 14501 23151
rect 14621 23150 14691 23151
rect 14041 23140 14910 23150
rect 14041 23132 14830 23140
rect 14041 23050 14050 23132
rect 14102 23050 14250 23132
rect 14302 23050 14440 23132
rect 14492 23050 14630 23132
rect 14682 23050 14830 23132
rect 14041 23040 14830 23050
rect 14900 23040 14910 23140
rect 15901 23090 15910 23172
rect 15962 23090 16100 23172
rect 16152 23090 16161 23172
rect 15901 23071 16161 23090
rect 15920 23070 16160 23071
rect 14041 23031 14910 23040
rect 14060 23030 14910 23031
rect 13648 23028 13802 23030
rect 16316 22170 16444 23410
rect 17213 22170 17283 22173
rect 17412 22170 17482 22171
rect 17603 22170 17673 22172
rect 16316 22163 17673 22170
rect 16316 22160 17220 22163
rect 16316 22049 16658 22160
rect 16711 22049 16839 22160
rect 16892 22049 17029 22160
rect 17082 22052 17220 22160
rect 17273 22162 17673 22163
rect 17273 22161 17610 22162
rect 17273 22052 17419 22161
rect 17082 22050 17419 22052
rect 17472 22051 17610 22161
rect 17663 22051 17673 22162
rect 17472 22050 17673 22051
rect 17082 22049 17673 22050
rect 16316 22042 17673 22049
rect 16650 22040 17660 22042
rect 18170 21356 18480 25024
rect 16840 21322 18481 21356
rect 15801 21310 15871 21311
rect 16001 21310 16071 21311
rect 15801 21292 16071 21310
rect 15801 21274 15810 21292
rect 13964 21271 15810 21274
rect 13951 21252 15810 21271
rect 13951 21170 13960 21252
rect 14012 21170 14150 21252
rect 14202 21170 14340 21252
rect 14392 21170 14530 21252
rect 14582 21170 14730 21252
rect 14782 21210 15810 21252
rect 15862 21210 16010 21292
rect 16062 21274 16071 21292
rect 16062 21210 16074 21274
rect 14782 21170 16074 21210
rect 12358 21112 12859 21158
rect 13951 21151 16074 21170
rect 13964 21146 16074 21151
rect 12358 20456 12405 21112
rect 12821 20903 12859 21112
rect 15615 20903 15745 21146
rect 16840 20932 16864 21322
rect 17006 20932 18481 21322
rect 12821 20731 15766 20903
rect 16840 20902 18481 20932
rect 12821 20456 12859 20731
rect 14540 20550 15490 20570
rect 14540 20490 14920 20550
rect 15460 20490 15490 20550
rect 14540 20470 15490 20490
rect 12358 20416 12859 20456
rect 14550 20020 14650 20470
rect 15615 20440 15745 20731
rect 14900 20430 15745 20440
rect 14900 20320 14910 20430
rect 14970 20320 15100 20430
rect 15160 20320 15300 20430
rect 15360 20320 15490 20430
rect 15550 20320 15745 20430
rect 14900 20310 15745 20320
rect 13010 19920 14650 20020
rect 15615 19965 15745 20310
rect 15615 19960 16175 19965
rect 15615 19950 16330 19960
rect 12531 17968 12811 17995
rect 12531 17700 12559 17968
rect 12791 17700 12811 17968
rect 12531 17677 12811 17700
rect 12640 17100 12940 17130
rect 12640 16860 12660 17100
rect 12910 17080 12940 17100
rect 13010 17080 13110 19920
rect 15615 19840 16070 19950
rect 16130 19840 16260 19950
rect 16320 19840 16330 19950
rect 15615 19835 16175 19840
rect 16060 19830 16140 19835
rect 16250 19830 16330 19840
rect 14810 19290 15460 19300
rect 14810 19180 14820 19290
rect 14880 19180 15010 19290
rect 15070 19180 15200 19290
rect 15260 19180 15390 19290
rect 15450 19180 15460 19290
rect 14810 19170 15460 19180
rect 15960 19280 16040 19290
rect 16160 19280 16240 19290
rect 15960 19170 15970 19280
rect 16030 19170 16170 19280
rect 16230 19260 17230 19280
rect 16230 19170 17040 19260
rect 17210 19170 17230 19260
rect 15960 19160 17230 19170
rect 16490 19120 16620 19130
rect 16490 19030 16500 19120
rect 16600 19030 16620 19120
rect 16490 19020 16620 19030
rect 16500 18050 16620 19020
rect 18200 19070 18590 19110
rect 18200 18985 18230 19070
rect 17725 18695 18230 18985
rect 17330 18050 17530 18060
rect 16500 18040 17530 18050
rect 16500 17940 16790 18040
rect 16870 17940 17350 18040
rect 16500 17930 17350 17940
rect 14642 17835 15187 17851
rect 14642 17833 15115 17835
rect 14642 17606 14654 17833
rect 14737 17606 15115 17833
rect 15175 17606 15187 17835
rect 17330 17740 17350 17930
rect 17510 17740 17530 18040
rect 17330 17720 17530 17740
rect 14642 17594 15187 17606
rect 17725 17570 18015 18695
rect 18200 18610 18230 18695
rect 18560 18985 18590 19070
rect 18560 18695 18635 18985
rect 18560 18610 18590 18695
rect 18200 18580 18590 18610
rect 16720 17566 17230 17570
rect 17270 17566 18020 17570
rect 16720 17530 18020 17566
rect 16720 17300 16760 17530
rect 16950 17300 18020 17530
rect 16720 17286 18020 17300
rect 16720 17280 17230 17286
rect 17270 17280 18020 17286
rect 18110 17283 18521 17306
rect 18110 17205 18146 17283
rect 12910 16980 13110 17080
rect 16741 17045 18146 17205
rect 12910 16860 12940 16980
rect 12640 16830 12940 16860
rect 16741 16714 16901 17045
rect 18110 17007 18146 17045
rect 18491 17007 18521 17283
rect 18110 16980 18521 17007
rect 12860 16694 16901 16714
rect 12860 16574 14156 16694
rect 14286 16692 16901 16694
rect 14286 16574 15456 16692
rect 12860 16566 15456 16574
rect 15515 16566 16901 16692
rect 12860 16554 16901 16566
rect 12490 16110 12770 16140
rect 12490 15790 12510 16110
rect 12750 16000 12770 16110
rect 12860 16000 13020 16554
rect 13506 16384 13602 16397
rect 13506 16289 13528 16384
rect 13592 16289 13602 16384
rect 13506 16279 13602 16289
rect 14486 16264 14646 16554
rect 15016 16484 15126 16494
rect 15016 16284 15026 16484
rect 15116 16284 15126 16484
rect 15016 16274 15126 16284
rect 14486 16234 14966 16264
rect 14486 16104 15196 16234
rect 12750 15840 13020 16000
rect 13119 16070 14305 16073
rect 13119 16004 14844 16070
rect 13119 15944 14752 16004
rect 14832 15944 14844 16004
rect 13119 15932 14844 15944
rect 13119 15851 14305 15932
rect 15036 15904 15196 16104
rect 14486 15894 15196 15904
rect 12750 15790 12770 15840
rect 12490 15770 12770 15790
rect 12512 14257 12732 14258
rect 13119 14257 13341 15851
rect 14486 15794 14502 15894
rect 14554 15794 14702 15894
rect 14754 15794 14892 15894
rect 14944 15794 15082 15894
rect 15134 15794 15196 15894
rect 17173 15934 17433 15944
rect 17173 15834 17182 15934
rect 17234 15834 17372 15934
rect 17424 15834 17433 15934
rect 17173 15824 17433 15834
rect 14486 15784 14646 15794
rect 14693 15784 14763 15794
rect 14883 15784 14953 15794
rect 15073 15784 15143 15794
rect 13507 15439 13602 15452
rect 13507 15320 13520 15439
rect 13589 15320 13602 15439
rect 13507 15307 13602 15320
rect 12512 14036 13341 14257
rect 12512 10620 12733 14036
rect 13119 14035 13341 14036
rect 17073 14054 17343 14064
rect 14413 14029 14483 14034
rect 14593 14029 14663 14034
rect 14783 14029 14853 14034
rect 14973 14029 15043 14034
rect 15163 14029 15233 14034
rect 14413 14024 15233 14029
rect 14413 13924 14422 14024
rect 14474 13924 14602 14024
rect 14654 13924 14792 14024
rect 14844 13924 14982 14024
rect 15034 13924 15172 14024
rect 15224 13924 15233 14024
rect 17073 13954 17082 14054
rect 17134 13954 17282 14054
rect 17334 13954 17343 14054
rect 17073 13944 17343 13954
rect 14413 13914 15233 13924
rect 14419 13911 15227 13914
rect 12862 13883 13120 13900
rect 12862 13871 13662 13883
rect 12862 13864 13668 13871
rect 12862 13803 13611 13864
rect 13663 13803 13668 13864
rect 12862 13794 13668 13803
rect 12862 13745 13662 13794
rect 12482 10608 12760 10620
rect 12862 10612 13120 13745
rect 14672 13071 14862 13911
rect 17132 13071 17332 13944
rect 13519 13070 17434 13071
rect 13519 13062 17446 13070
rect 13508 13058 17446 13062
rect 13508 13057 14216 13058
rect 13508 13055 14042 13057
rect 13508 13052 13685 13055
rect 13508 12960 13512 13052
rect 13566 12966 13685 13052
rect 13737 13052 14042 13055
rect 13737 12966 13860 13052
rect 13566 12960 13860 12966
rect 13914 12968 14042 13052
rect 14094 12968 14216 13057
rect 13914 12966 14216 12968
rect 14270 13057 14747 13058
rect 14270 12968 14395 13057
rect 14447 13056 14747 13057
rect 14447 12968 14566 13056
rect 14270 12966 14566 12968
rect 13914 12964 14566 12966
rect 14620 12969 14747 13056
rect 14799 13057 15274 13058
rect 14799 13056 15098 13057
rect 14799 12969 14920 13056
rect 14620 12964 14920 12969
rect 14974 12968 15098 13056
rect 15150 12968 15274 13057
rect 14974 12966 15274 12968
rect 15328 13052 15626 13058
rect 15328 12966 15450 13052
rect 14974 12964 15450 12966
rect 13914 12963 15450 12964
rect 15502 12966 15626 13052
rect 15680 13057 17446 13058
rect 15680 13056 16858 13057
rect 15680 13054 16680 13056
rect 15680 13052 15976 13054
rect 15680 12966 15803 13052
rect 15502 12963 15803 12966
rect 15855 12963 15976 13052
rect 13914 12962 15976 12963
rect 16030 13052 16330 13054
rect 16030 12963 16155 13052
rect 16207 12963 16330 13052
rect 16030 12962 16330 12963
rect 16384 13051 16680 13054
rect 16384 12962 16509 13051
rect 16561 12964 16680 13051
rect 16734 12968 16858 13056
rect 16910 13056 17388 13057
rect 16910 12968 17034 13056
rect 16734 12964 17034 12968
rect 17088 13052 17388 13056
rect 17088 12964 17211 13052
rect 16561 12963 17211 12964
rect 17263 12968 17388 13052
rect 17440 12968 17446 13057
rect 17263 12963 17446 12968
rect 16561 12962 17446 12963
rect 13914 12960 17446 12962
rect 13508 12956 17446 12960
rect 13508 12950 13570 12956
rect 13678 12954 13743 12956
rect 13856 12950 13918 12956
rect 14562 12954 14624 12956
rect 14672 12954 14862 12956
rect 14916 12954 14978 12956
rect 15443 12951 15508 12956
rect 15796 12951 15861 12956
rect 15972 12952 16034 12956
rect 16148 12951 16213 12956
rect 16326 12952 16388 12956
rect 16502 12950 16567 12956
rect 16676 12954 16738 12956
rect 17030 12954 17092 12956
rect 17204 12951 17269 12956
rect 17262 10624 17568 10784
rect 12482 10354 12496 10608
rect 12738 10354 12760 10608
rect 12856 10598 13126 10612
rect 12856 10366 12868 10598
rect 13112 10366 13126 10598
rect 12856 10356 13126 10366
rect 17262 10372 17276 10624
rect 17542 10372 17568 10624
rect 17262 10356 17568 10372
rect 17792 10640 18052 10712
rect 17792 10380 17806 10640
rect 18034 10380 18052 10640
rect 17792 10366 18052 10380
rect 12868 10354 13126 10356
rect 12482 10342 12760 10354
rect 4162 8388 4218 9718
rect 5576 8388 5612 9718
rect 4162 8324 5612 8388
rect 25230 9698 26614 25642
rect 25230 8378 25266 9698
rect 26538 8378 26614 9698
rect 25230 8342 26614 8378
rect 2168 6346 2324 7480
rect 3678 6346 3820 7480
rect 2168 6246 3820 6346
rect 27052 7470 28704 27758
rect 27052 6336 27174 7470
rect 28528 6336 28704 7470
rect 27052 6246 28704 6336
<< via2 >>
rect 12340 24874 12564 25304
rect 17844 25110 18020 25332
rect 18192 25024 18456 25302
rect 15272 23364 15414 23612
rect 12405 20456 12821 21112
rect 12559 17700 12791 17968
rect 12660 16860 12910 17100
rect 17350 17740 17510 18040
rect 18230 18610 18560 19070
rect 18146 17007 18491 17283
rect 12510 15790 12750 16110
rect 13528 16289 13592 16384
rect 15026 16284 15116 16484
rect 13520 15320 13589 15439
rect 12496 10354 12738 10608
rect 12868 10366 13112 10598
rect 17276 10372 17542 10624
rect 17806 10380 18034 10640
<< metal3 >>
rect 17830 25332 18030 25342
rect 11908 24682 12188 25328
rect 12322 25304 12584 25328
rect 12322 24874 12340 25304
rect 12564 24874 12584 25304
rect 17830 25110 17844 25332
rect 18020 25110 18030 25332
rect 17830 25096 18030 25110
rect 18168 25302 18478 25326
rect 18168 25024 18192 25302
rect 18456 25024 18478 25302
rect 18168 25006 18478 25024
rect 12322 24852 12584 24874
rect 11908 24402 12448 24682
rect 12168 23630 12448 24402
rect 12168 23612 15432 23630
rect 12168 23364 15272 23612
rect 15414 23364 15432 23612
rect 12168 23350 15432 23364
rect 12358 21112 12859 21158
rect 12358 20456 12405 21112
rect 12821 20456 12859 21112
rect 12358 20416 12859 20456
rect 18200 19070 18590 19110
rect 18200 18610 18230 19070
rect 18560 18610 18590 19070
rect 18200 18580 18590 18610
rect 17330 18040 17530 18060
rect 12531 17968 12811 17995
rect 12531 17700 12559 17968
rect 12791 17700 12811 17968
rect 17330 17740 17350 18040
rect 17510 17740 17530 18040
rect 17330 17720 17530 17740
rect 12531 17677 12811 17700
rect 18110 17283 18521 17306
rect 12640 17100 12940 17130
rect 12640 16860 12660 17100
rect 12910 16860 12940 17100
rect 18110 17007 18146 17283
rect 18491 17007 18521 17283
rect 18110 16980 18521 17007
rect 12640 16830 12940 16860
rect 18316 16584 18586 16614
rect 18316 16499 18336 16584
rect 15015 16484 18336 16499
rect 13507 16384 13602 16396
rect 13507 16289 13528 16384
rect 13592 16289 13602 16384
rect 12490 16110 12770 16140
rect 12490 15790 12510 16110
rect 12750 15790 12770 16110
rect 12490 15770 12770 15790
rect 13507 15439 13602 16289
rect 15015 16288 15026 16484
rect 15016 16284 15026 16288
rect 15116 16288 18336 16484
rect 15116 16284 15126 16288
rect 15016 16274 15126 16284
rect 18316 16254 18336 16288
rect 18566 16254 18586 16584
rect 18316 16224 18586 16254
rect 13507 15320 13520 15439
rect 13589 15320 13602 15439
rect 13507 15307 13602 15320
rect 17262 10624 17568 10784
rect 12482 10608 12760 10620
rect 12482 10354 12496 10608
rect 12738 10354 12760 10608
rect 12862 10598 13120 10604
rect 12862 10366 12868 10598
rect 13112 10366 13120 10598
rect 12862 10360 13120 10366
rect 17262 10372 17276 10624
rect 17542 10372 17568 10624
rect 17262 10356 17568 10372
rect 17792 10640 18052 10712
rect 17792 10380 17806 10640
rect 18034 10380 18052 10640
rect 17792 10366 18052 10380
rect 12482 10342 12760 10354
<< via3 >>
rect 12405 20456 12821 21112
rect 18230 18610 18560 19070
rect 12559 17700 12791 17968
rect 17350 17740 17510 18040
rect 12660 16860 12910 17100
rect 18146 17007 18491 17283
rect 12510 15790 12750 16110
rect 18336 16254 18566 16584
<< metal4 >>
rect 5947 17996 12147 24400
rect 12358 21112 12859 21158
rect 12358 20456 12405 21112
rect 12821 20456 12859 21112
rect 12358 20416 12859 20456
rect 18200 19070 18590 19110
rect 18200 18610 18230 19070
rect 18560 18610 18590 19070
rect 18200 18580 18590 18610
rect 18861 18060 25061 24454
rect 17330 18040 25061 18060
rect 5947 17968 12813 17996
rect 5947 17954 12559 17968
rect 5947 17718 5988 17954
rect 12106 17718 12559 17954
rect 5947 17700 12559 17718
rect 12791 17700 12813 17968
rect 17330 17740 17350 18040
rect 17510 18008 25061 18040
rect 17510 17772 18902 18008
rect 25020 17772 25061 18008
rect 17510 17752 25061 17772
rect 17510 17740 19240 17752
rect 17330 17720 19240 17740
rect 5947 17698 12813 17700
rect 11905 17677 12813 17698
rect 18110 17283 19228 17305
rect 5991 17130 12191 17132
rect 5991 17112 12940 17130
rect 5991 16876 6032 17112
rect 12150 17100 12940 17112
rect 12150 16876 12660 17100
rect 5991 16860 12660 16876
rect 12910 16860 12940 17100
rect 18110 17007 18146 17283
rect 18491 17282 19228 17283
rect 18491 17262 25060 17282
rect 18491 17026 18901 17262
rect 25019 17026 25060 17262
rect 18491 17007 25060 17026
rect 18110 16980 25060 17007
rect 5991 16830 12940 16860
rect 5991 10430 12191 16830
rect 18316 16585 18586 16614
rect 18316 16252 18332 16585
rect 18572 16252 18586 16585
rect 18316 16224 18586 16252
rect 12490 16110 12770 16140
rect 12490 15790 12510 16110
rect 12750 15790 12770 16110
rect 12490 15770 12770 15790
rect 18860 10580 25060 16980
<< via4 >>
rect 12405 20456 12821 21112
rect 18230 18610 18560 19070
rect 5988 17718 12106 17954
rect 18902 17772 25020 18008
rect 6032 16876 12150 17112
rect 18901 17026 25019 17262
rect 18332 16584 18572 16585
rect 18332 16254 18336 16584
rect 18336 16254 18566 16584
rect 18566 16254 18572 16584
rect 18332 16252 18572 16254
rect 12510 15790 12750 16110
<< mimcap2 >>
rect 18961 24314 24961 24354
rect 6047 24260 12047 24300
rect 6047 18340 6087 24260
rect 12007 18340 12047 24260
rect 18961 18394 19001 24314
rect 24921 18394 24961 24314
rect 18961 18354 24961 18394
rect 6047 18300 12047 18340
rect 18960 16640 24960 16680
rect 6091 16490 12091 16530
rect 6091 10570 6131 16490
rect 12051 10570 12091 16490
rect 18960 10720 19000 16640
rect 24920 10720 24960 16640
rect 18960 10680 24960 10720
rect 6091 10530 12091 10570
<< mimcap2contact >>
rect 6087 18340 12007 24260
rect 19001 18394 24921 24314
rect 6131 10570 12051 16490
rect 19000 10720 24920 16640
<< metal5 >>
rect 18977 24314 24945 24338
rect 6063 24260 12031 24284
rect 6063 18340 6087 24260
rect 12007 21154 12031 24260
rect 12007 21112 12857 21154
rect 12007 20456 12405 21112
rect 12821 20456 12857 21112
rect 12007 20418 12857 20456
rect 12007 18340 12031 20418
rect 18977 19110 19001 24314
rect 18200 19070 19001 19110
rect 18200 18610 18230 19070
rect 18560 18610 19001 19070
rect 18200 18580 19001 18610
rect 18977 18394 19001 18580
rect 24921 18394 24945 24314
rect 18977 18370 24945 18394
rect 6063 18316 12031 18340
rect 18860 18008 25062 18050
rect 5946 17954 12148 17996
rect 5946 17718 5988 17954
rect 12106 17718 12148 17954
rect 18860 17772 18902 18008
rect 25020 17772 25062 18008
rect 18860 17730 25062 17772
rect 5946 17676 12148 17718
rect 18859 17262 25061 17304
rect 5990 17112 12192 17154
rect 5990 16876 6032 17112
rect 12150 16876 12192 17112
rect 18859 17026 18901 17262
rect 25019 17026 25061 17262
rect 18859 16984 25061 17026
rect 5990 16834 12192 16876
rect 18976 16640 24944 16664
rect 18976 16614 19000 16640
rect 18281 16585 19000 16614
rect 6107 16490 12075 16514
rect 6107 10570 6131 16490
rect 12051 16160 12075 16490
rect 18281 16252 18332 16585
rect 18572 16252 19000 16585
rect 18281 16224 19000 16252
rect 12051 16110 12800 16160
rect 12051 15790 12510 16110
rect 12750 15790 12800 16110
rect 12051 15750 12800 15790
rect 12051 10570 12075 15750
rect 18976 10720 19000 16224
rect 24920 10720 24944 16640
rect 18976 10696 24944 10720
rect 6107 10546 12075 10570
<< res0p35 >>
rect 13476 24544 16480 24618
rect 13506 23864 14310 23938
rect 13484 21536 13558 21640
rect 15304 21556 15378 22800
rect 16784 19316 16858 20920
rect 14640 17320 14714 17424
rect 15860 17320 15934 17424
rect 16252 17321 16326 18125
rect 17394 17936 17468 20940
rect 16146 14290 16220 15534
<< res0p69 >>
rect 13742 19590 13884 19732
rect 13742 19204 13884 19346
rect 13742 18818 13884 18960
rect 13742 18432 13884 18574
rect 13742 18046 13884 18188
rect 13742 17660 13884 17802
rect 13742 17274 13884 17416
rect 13742 16888 13884 17030
<< labels >>
flabel metal3 12000 25086 12000 25086 0 FreeSans 1280 90 0 0 VB0_6
port 10 nsew
flabel via2 12442 25032 12442 25032 0 FreeSans 1280 90 0 0 VSI2
port 9 nsew
flabel locali 14542 25052 14542 25052 0 FreeSans 1280 90 0 0 VDD
port 6 nsew
flabel via2 17928 25256 17928 25256 0 FreeSans 1280 90 0 0 VOUT
port 11 nsew
flabel via2 18282 25126 18282 25126 0 FreeSans 1280 90 0 0 VB0_9
port 8 nsew
flabel locali 15294 10468 15294 10468 0 FreeSans 1280 90 0 0 VSS
port 2 nsew
flabel via2 17420 10482 17420 10482 0 FreeSans 1280 90 0 0 VSI1
port 4 nsew
flabel via2 17906 10532 17906 10532 0 FreeSans 1280 90 0 0 VB1_5
port 7 nsew
flabel via2 13002 10468 13002 10468 0 FreeSans 1280 90 0 0 VB0_75
port 3 nsew
flabel via2 12582 10524 12582 10524 0 FreeSans 1280 90 0 0 VB1_4
port 5 nsew
flabel metal1 13510 10494 13518 10494 0 FreeSans 1600 90 0 0 VRF
port 1 nsew
<< end >>
