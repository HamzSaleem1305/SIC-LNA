magic
tech sky130A
magscale 1 2
timestamp 1666356932
<< error_p >>
rect -893 1120 -835 1126
rect -701 1120 -643 1126
rect -509 1120 -451 1126
rect -317 1120 -259 1126
rect -125 1120 -67 1126
rect 67 1120 125 1126
rect 259 1120 317 1126
rect 451 1120 509 1126
rect 643 1120 701 1126
rect 835 1120 893 1126
rect -893 1086 -881 1120
rect -701 1086 -689 1120
rect -509 1086 -497 1120
rect -317 1086 -305 1120
rect -125 1086 -113 1120
rect 67 1086 79 1120
rect 259 1086 271 1120
rect 451 1086 463 1120
rect 643 1086 655 1120
rect 835 1086 847 1120
rect -893 1080 -835 1086
rect -701 1080 -643 1086
rect -509 1080 -451 1086
rect -317 1080 -259 1086
rect -125 1080 -67 1086
rect 67 1080 125 1086
rect 259 1080 317 1086
rect 451 1080 509 1086
rect 643 1080 701 1086
rect 835 1080 893 1086
rect -989 -1086 -931 -1080
rect -797 -1086 -739 -1080
rect -605 -1086 -547 -1080
rect -413 -1086 -355 -1080
rect -221 -1086 -163 -1080
rect -29 -1086 29 -1080
rect 163 -1086 221 -1080
rect 355 -1086 413 -1080
rect 547 -1086 605 -1080
rect 739 -1086 797 -1080
rect 931 -1086 989 -1080
rect -989 -1120 -977 -1086
rect -797 -1120 -785 -1086
rect -605 -1120 -593 -1086
rect -413 -1120 -401 -1086
rect -221 -1120 -209 -1086
rect -29 -1120 -17 -1086
rect 163 -1120 175 -1086
rect 355 -1120 367 -1086
rect 547 -1120 559 -1086
rect 739 -1120 751 -1086
rect 931 -1120 943 -1086
rect -989 -1126 -931 -1120
rect -797 -1126 -739 -1120
rect -605 -1126 -547 -1120
rect -413 -1126 -355 -1120
rect -221 -1126 -163 -1120
rect -29 -1126 29 -1120
rect 163 -1126 221 -1120
rect 355 -1126 413 -1120
rect 547 -1126 605 -1120
rect 739 -1126 797 -1120
rect 931 -1126 989 -1120
<< pwell >>
rect -1175 -1258 1175 1258
<< nmoslvt >>
rect -975 -1048 -945 1048
rect -879 -1048 -849 1048
rect -783 -1048 -753 1048
rect -687 -1048 -657 1048
rect -591 -1048 -561 1048
rect -495 -1048 -465 1048
rect -399 -1048 -369 1048
rect -303 -1048 -273 1048
rect -207 -1048 -177 1048
rect -111 -1048 -81 1048
rect -15 -1048 15 1048
rect 81 -1048 111 1048
rect 177 -1048 207 1048
rect 273 -1048 303 1048
rect 369 -1048 399 1048
rect 465 -1048 495 1048
rect 561 -1048 591 1048
rect 657 -1048 687 1048
rect 753 -1048 783 1048
rect 849 -1048 879 1048
rect 945 -1048 975 1048
<< ndiff >>
rect -1037 1036 -975 1048
rect -1037 -1036 -1025 1036
rect -991 -1036 -975 1036
rect -1037 -1048 -975 -1036
rect -945 1036 -879 1048
rect -945 -1036 -929 1036
rect -895 -1036 -879 1036
rect -945 -1048 -879 -1036
rect -849 1036 -783 1048
rect -849 -1036 -833 1036
rect -799 -1036 -783 1036
rect -849 -1048 -783 -1036
rect -753 1036 -687 1048
rect -753 -1036 -737 1036
rect -703 -1036 -687 1036
rect -753 -1048 -687 -1036
rect -657 1036 -591 1048
rect -657 -1036 -641 1036
rect -607 -1036 -591 1036
rect -657 -1048 -591 -1036
rect -561 1036 -495 1048
rect -561 -1036 -545 1036
rect -511 -1036 -495 1036
rect -561 -1048 -495 -1036
rect -465 1036 -399 1048
rect -465 -1036 -449 1036
rect -415 -1036 -399 1036
rect -465 -1048 -399 -1036
rect -369 1036 -303 1048
rect -369 -1036 -353 1036
rect -319 -1036 -303 1036
rect -369 -1048 -303 -1036
rect -273 1036 -207 1048
rect -273 -1036 -257 1036
rect -223 -1036 -207 1036
rect -273 -1048 -207 -1036
rect -177 1036 -111 1048
rect -177 -1036 -161 1036
rect -127 -1036 -111 1036
rect -177 -1048 -111 -1036
rect -81 1036 -15 1048
rect -81 -1036 -65 1036
rect -31 -1036 -15 1036
rect -81 -1048 -15 -1036
rect 15 1036 81 1048
rect 15 -1036 31 1036
rect 65 -1036 81 1036
rect 15 -1048 81 -1036
rect 111 1036 177 1048
rect 111 -1036 127 1036
rect 161 -1036 177 1036
rect 111 -1048 177 -1036
rect 207 1036 273 1048
rect 207 -1036 223 1036
rect 257 -1036 273 1036
rect 207 -1048 273 -1036
rect 303 1036 369 1048
rect 303 -1036 319 1036
rect 353 -1036 369 1036
rect 303 -1048 369 -1036
rect 399 1036 465 1048
rect 399 -1036 415 1036
rect 449 -1036 465 1036
rect 399 -1048 465 -1036
rect 495 1036 561 1048
rect 495 -1036 511 1036
rect 545 -1036 561 1036
rect 495 -1048 561 -1036
rect 591 1036 657 1048
rect 591 -1036 607 1036
rect 641 -1036 657 1036
rect 591 -1048 657 -1036
rect 687 1036 753 1048
rect 687 -1036 703 1036
rect 737 -1036 753 1036
rect 687 -1048 753 -1036
rect 783 1036 849 1048
rect 783 -1036 799 1036
rect 833 -1036 849 1036
rect 783 -1048 849 -1036
rect 879 1036 945 1048
rect 879 -1036 895 1036
rect 929 -1036 945 1036
rect 879 -1048 945 -1036
rect 975 1036 1037 1048
rect 975 -1036 991 1036
rect 1025 -1036 1037 1036
rect 975 -1048 1037 -1036
<< ndiffc >>
rect -1025 -1036 -991 1036
rect -929 -1036 -895 1036
rect -833 -1036 -799 1036
rect -737 -1036 -703 1036
rect -641 -1036 -607 1036
rect -545 -1036 -511 1036
rect -449 -1036 -415 1036
rect -353 -1036 -319 1036
rect -257 -1036 -223 1036
rect -161 -1036 -127 1036
rect -65 -1036 -31 1036
rect 31 -1036 65 1036
rect 127 -1036 161 1036
rect 223 -1036 257 1036
rect 319 -1036 353 1036
rect 415 -1036 449 1036
rect 511 -1036 545 1036
rect 607 -1036 641 1036
rect 703 -1036 737 1036
rect 799 -1036 833 1036
rect 895 -1036 929 1036
rect 991 -1036 1025 1036
<< psubdiff >>
rect -1139 1188 -1043 1222
rect 1043 1188 1139 1222
rect -1139 1126 -1105 1188
rect 1105 1126 1139 1188
rect -1139 -1188 -1105 -1126
rect 1105 -1188 1139 -1126
rect -1139 -1222 -1043 -1188
rect 1043 -1222 1139 -1188
<< psubdiffcont >>
rect -1043 1188 1043 1222
rect -1139 -1126 -1105 1126
rect 1105 -1126 1139 1126
rect -1043 -1222 1043 -1188
<< poly >>
rect -897 1120 -831 1136
rect -897 1086 -881 1120
rect -847 1086 -831 1120
rect -975 1048 -945 1074
rect -897 1070 -831 1086
rect -705 1120 -639 1136
rect -705 1086 -689 1120
rect -655 1086 -639 1120
rect -879 1048 -849 1070
rect -783 1048 -753 1074
rect -705 1070 -639 1086
rect -513 1120 -447 1136
rect -513 1086 -497 1120
rect -463 1086 -447 1120
rect -687 1048 -657 1070
rect -591 1048 -561 1074
rect -513 1070 -447 1086
rect -321 1120 -255 1136
rect -321 1086 -305 1120
rect -271 1086 -255 1120
rect -495 1048 -465 1070
rect -399 1048 -369 1074
rect -321 1070 -255 1086
rect -129 1120 -63 1136
rect -129 1086 -113 1120
rect -79 1086 -63 1120
rect -303 1048 -273 1070
rect -207 1048 -177 1074
rect -129 1070 -63 1086
rect 63 1120 129 1136
rect 63 1086 79 1120
rect 113 1086 129 1120
rect -111 1048 -81 1070
rect -15 1048 15 1074
rect 63 1070 129 1086
rect 255 1120 321 1136
rect 255 1086 271 1120
rect 305 1086 321 1120
rect 81 1048 111 1070
rect 177 1048 207 1074
rect 255 1070 321 1086
rect 447 1120 513 1136
rect 447 1086 463 1120
rect 497 1086 513 1120
rect 273 1048 303 1070
rect 369 1048 399 1074
rect 447 1070 513 1086
rect 639 1120 705 1136
rect 639 1086 655 1120
rect 689 1086 705 1120
rect 465 1048 495 1070
rect 561 1048 591 1074
rect 639 1070 705 1086
rect 831 1120 897 1136
rect 831 1086 847 1120
rect 881 1086 897 1120
rect 657 1048 687 1070
rect 753 1048 783 1074
rect 831 1070 897 1086
rect 849 1048 879 1070
rect 945 1048 975 1074
rect -975 -1070 -945 -1048
rect -993 -1086 -927 -1070
rect -879 -1074 -849 -1048
rect -783 -1070 -753 -1048
rect -993 -1120 -977 -1086
rect -943 -1120 -927 -1086
rect -993 -1136 -927 -1120
rect -801 -1086 -735 -1070
rect -687 -1074 -657 -1048
rect -591 -1070 -561 -1048
rect -801 -1120 -785 -1086
rect -751 -1120 -735 -1086
rect -801 -1136 -735 -1120
rect -609 -1086 -543 -1070
rect -495 -1074 -465 -1048
rect -399 -1070 -369 -1048
rect -609 -1120 -593 -1086
rect -559 -1120 -543 -1086
rect -609 -1136 -543 -1120
rect -417 -1086 -351 -1070
rect -303 -1074 -273 -1048
rect -207 -1070 -177 -1048
rect -417 -1120 -401 -1086
rect -367 -1120 -351 -1086
rect -417 -1136 -351 -1120
rect -225 -1086 -159 -1070
rect -111 -1074 -81 -1048
rect -15 -1070 15 -1048
rect -225 -1120 -209 -1086
rect -175 -1120 -159 -1086
rect -225 -1136 -159 -1120
rect -33 -1086 33 -1070
rect 81 -1074 111 -1048
rect 177 -1070 207 -1048
rect -33 -1120 -17 -1086
rect 17 -1120 33 -1086
rect -33 -1136 33 -1120
rect 159 -1086 225 -1070
rect 273 -1074 303 -1048
rect 369 -1070 399 -1048
rect 159 -1120 175 -1086
rect 209 -1120 225 -1086
rect 159 -1136 225 -1120
rect 351 -1086 417 -1070
rect 465 -1074 495 -1048
rect 561 -1070 591 -1048
rect 351 -1120 367 -1086
rect 401 -1120 417 -1086
rect 351 -1136 417 -1120
rect 543 -1086 609 -1070
rect 657 -1074 687 -1048
rect 753 -1070 783 -1048
rect 543 -1120 559 -1086
rect 593 -1120 609 -1086
rect 543 -1136 609 -1120
rect 735 -1086 801 -1070
rect 849 -1074 879 -1048
rect 945 -1070 975 -1048
rect 735 -1120 751 -1086
rect 785 -1120 801 -1086
rect 735 -1136 801 -1120
rect 927 -1086 993 -1070
rect 927 -1120 943 -1086
rect 977 -1120 993 -1086
rect 927 -1136 993 -1120
<< polycont >>
rect -881 1086 -847 1120
rect -689 1086 -655 1120
rect -497 1086 -463 1120
rect -305 1086 -271 1120
rect -113 1086 -79 1120
rect 79 1086 113 1120
rect 271 1086 305 1120
rect 463 1086 497 1120
rect 655 1086 689 1120
rect 847 1086 881 1120
rect -977 -1120 -943 -1086
rect -785 -1120 -751 -1086
rect -593 -1120 -559 -1086
rect -401 -1120 -367 -1086
rect -209 -1120 -175 -1086
rect -17 -1120 17 -1086
rect 175 -1120 209 -1086
rect 367 -1120 401 -1086
rect 559 -1120 593 -1086
rect 751 -1120 785 -1086
rect 943 -1120 977 -1086
<< locali >>
rect -1139 1188 -1043 1222
rect 1043 1188 1139 1222
rect -1139 1126 -1105 1188
rect 1105 1126 1139 1188
rect -897 1086 -881 1120
rect -847 1086 -831 1120
rect -705 1086 -689 1120
rect -655 1086 -639 1120
rect -513 1086 -497 1120
rect -463 1086 -447 1120
rect -321 1086 -305 1120
rect -271 1086 -255 1120
rect -129 1086 -113 1120
rect -79 1086 -63 1120
rect 63 1086 79 1120
rect 113 1086 129 1120
rect 255 1086 271 1120
rect 305 1086 321 1120
rect 447 1086 463 1120
rect 497 1086 513 1120
rect 639 1086 655 1120
rect 689 1086 705 1120
rect 831 1086 847 1120
rect 881 1086 897 1120
rect -1025 1036 -991 1052
rect -1025 -1052 -991 -1036
rect -929 1036 -895 1052
rect -929 -1052 -895 -1036
rect -833 1036 -799 1052
rect -833 -1052 -799 -1036
rect -737 1036 -703 1052
rect -737 -1052 -703 -1036
rect -641 1036 -607 1052
rect -641 -1052 -607 -1036
rect -545 1036 -511 1052
rect -545 -1052 -511 -1036
rect -449 1036 -415 1052
rect -449 -1052 -415 -1036
rect -353 1036 -319 1052
rect -353 -1052 -319 -1036
rect -257 1036 -223 1052
rect -257 -1052 -223 -1036
rect -161 1036 -127 1052
rect -161 -1052 -127 -1036
rect -65 1036 -31 1052
rect -65 -1052 -31 -1036
rect 31 1036 65 1052
rect 31 -1052 65 -1036
rect 127 1036 161 1052
rect 127 -1052 161 -1036
rect 223 1036 257 1052
rect 223 -1052 257 -1036
rect 319 1036 353 1052
rect 319 -1052 353 -1036
rect 415 1036 449 1052
rect 415 -1052 449 -1036
rect 511 1036 545 1052
rect 511 -1052 545 -1036
rect 607 1036 641 1052
rect 607 -1052 641 -1036
rect 703 1036 737 1052
rect 703 -1052 737 -1036
rect 799 1036 833 1052
rect 799 -1052 833 -1036
rect 895 1036 929 1052
rect 895 -1052 929 -1036
rect 991 1036 1025 1052
rect 991 -1052 1025 -1036
rect -993 -1120 -977 -1086
rect -943 -1120 -927 -1086
rect -801 -1120 -785 -1086
rect -751 -1120 -735 -1086
rect -609 -1120 -593 -1086
rect -559 -1120 -543 -1086
rect -417 -1120 -401 -1086
rect -367 -1120 -351 -1086
rect -225 -1120 -209 -1086
rect -175 -1120 -159 -1086
rect -33 -1120 -17 -1086
rect 17 -1120 33 -1086
rect 159 -1120 175 -1086
rect 209 -1120 225 -1086
rect 351 -1120 367 -1086
rect 401 -1120 417 -1086
rect 543 -1120 559 -1086
rect 593 -1120 609 -1086
rect 735 -1120 751 -1086
rect 785 -1120 801 -1086
rect 927 -1120 943 -1086
rect 977 -1120 993 -1086
rect -1139 -1188 -1105 -1126
rect 1105 -1188 1139 -1126
rect -1139 -1222 -1043 -1188
rect 1043 -1222 1139 -1188
<< viali >>
rect -881 1086 -847 1120
rect -689 1086 -655 1120
rect -497 1086 -463 1120
rect -305 1086 -271 1120
rect -113 1086 -79 1120
rect 79 1086 113 1120
rect 271 1086 305 1120
rect 463 1086 497 1120
rect 655 1086 689 1120
rect 847 1086 881 1120
rect -1025 -1036 -991 1036
rect -929 -1036 -895 1036
rect -833 -1036 -799 1036
rect -737 -1036 -703 1036
rect -641 -1036 -607 1036
rect -545 -1036 -511 1036
rect -449 -1036 -415 1036
rect -353 -1036 -319 1036
rect -257 -1036 -223 1036
rect -161 -1036 -127 1036
rect -65 -1036 -31 1036
rect 31 -1036 65 1036
rect 127 -1036 161 1036
rect 223 -1036 257 1036
rect 319 -1036 353 1036
rect 415 -1036 449 1036
rect 511 -1036 545 1036
rect 607 -1036 641 1036
rect 703 -1036 737 1036
rect 799 -1036 833 1036
rect 895 -1036 929 1036
rect 991 -1036 1025 1036
rect -977 -1120 -943 -1086
rect -785 -1120 -751 -1086
rect -593 -1120 -559 -1086
rect -401 -1120 -367 -1086
rect -209 -1120 -175 -1086
rect -17 -1120 17 -1086
rect 175 -1120 209 -1086
rect 367 -1120 401 -1086
rect 559 -1120 593 -1086
rect 751 -1120 785 -1086
rect 943 -1120 977 -1086
<< metal1 >>
rect -893 1120 -835 1126
rect -893 1086 -881 1120
rect -847 1086 -835 1120
rect -893 1080 -835 1086
rect -701 1120 -643 1126
rect -701 1086 -689 1120
rect -655 1086 -643 1120
rect -701 1080 -643 1086
rect -509 1120 -451 1126
rect -509 1086 -497 1120
rect -463 1086 -451 1120
rect -509 1080 -451 1086
rect -317 1120 -259 1126
rect -317 1086 -305 1120
rect -271 1086 -259 1120
rect -317 1080 -259 1086
rect -125 1120 -67 1126
rect -125 1086 -113 1120
rect -79 1086 -67 1120
rect -125 1080 -67 1086
rect 67 1120 125 1126
rect 67 1086 79 1120
rect 113 1086 125 1120
rect 67 1080 125 1086
rect 259 1120 317 1126
rect 259 1086 271 1120
rect 305 1086 317 1120
rect 259 1080 317 1086
rect 451 1120 509 1126
rect 451 1086 463 1120
rect 497 1086 509 1120
rect 451 1080 509 1086
rect 643 1120 701 1126
rect 643 1086 655 1120
rect 689 1086 701 1120
rect 643 1080 701 1086
rect 835 1120 893 1126
rect 835 1086 847 1120
rect 881 1086 893 1120
rect 835 1080 893 1086
rect -1031 1036 -985 1048
rect -1031 -1036 -1025 1036
rect -991 -1036 -985 1036
rect -1031 -1048 -985 -1036
rect -935 1036 -889 1048
rect -935 -1036 -929 1036
rect -895 -1036 -889 1036
rect -935 -1048 -889 -1036
rect -839 1036 -793 1048
rect -839 -1036 -833 1036
rect -799 -1036 -793 1036
rect -839 -1048 -793 -1036
rect -743 1036 -697 1048
rect -743 -1036 -737 1036
rect -703 -1036 -697 1036
rect -743 -1048 -697 -1036
rect -647 1036 -601 1048
rect -647 -1036 -641 1036
rect -607 -1036 -601 1036
rect -647 -1048 -601 -1036
rect -551 1036 -505 1048
rect -551 -1036 -545 1036
rect -511 -1036 -505 1036
rect -551 -1048 -505 -1036
rect -455 1036 -409 1048
rect -455 -1036 -449 1036
rect -415 -1036 -409 1036
rect -455 -1048 -409 -1036
rect -359 1036 -313 1048
rect -359 -1036 -353 1036
rect -319 -1036 -313 1036
rect -359 -1048 -313 -1036
rect -263 1036 -217 1048
rect -263 -1036 -257 1036
rect -223 -1036 -217 1036
rect -263 -1048 -217 -1036
rect -167 1036 -121 1048
rect -167 -1036 -161 1036
rect -127 -1036 -121 1036
rect -167 -1048 -121 -1036
rect -71 1036 -25 1048
rect -71 -1036 -65 1036
rect -31 -1036 -25 1036
rect -71 -1048 -25 -1036
rect 25 1036 71 1048
rect 25 -1036 31 1036
rect 65 -1036 71 1036
rect 25 -1048 71 -1036
rect 121 1036 167 1048
rect 121 -1036 127 1036
rect 161 -1036 167 1036
rect 121 -1048 167 -1036
rect 217 1036 263 1048
rect 217 -1036 223 1036
rect 257 -1036 263 1036
rect 217 -1048 263 -1036
rect 313 1036 359 1048
rect 313 -1036 319 1036
rect 353 -1036 359 1036
rect 313 -1048 359 -1036
rect 409 1036 455 1048
rect 409 -1036 415 1036
rect 449 -1036 455 1036
rect 409 -1048 455 -1036
rect 505 1036 551 1048
rect 505 -1036 511 1036
rect 545 -1036 551 1036
rect 505 -1048 551 -1036
rect 601 1036 647 1048
rect 601 -1036 607 1036
rect 641 -1036 647 1036
rect 601 -1048 647 -1036
rect 697 1036 743 1048
rect 697 -1036 703 1036
rect 737 -1036 743 1036
rect 697 -1048 743 -1036
rect 793 1036 839 1048
rect 793 -1036 799 1036
rect 833 -1036 839 1036
rect 793 -1048 839 -1036
rect 889 1036 935 1048
rect 889 -1036 895 1036
rect 929 -1036 935 1036
rect 889 -1048 935 -1036
rect 985 1036 1031 1048
rect 985 -1036 991 1036
rect 1025 -1036 1031 1036
rect 985 -1048 1031 -1036
rect -989 -1086 -931 -1080
rect -989 -1120 -977 -1086
rect -943 -1120 -931 -1086
rect -989 -1126 -931 -1120
rect -797 -1086 -739 -1080
rect -797 -1120 -785 -1086
rect -751 -1120 -739 -1086
rect -797 -1126 -739 -1120
rect -605 -1086 -547 -1080
rect -605 -1120 -593 -1086
rect -559 -1120 -547 -1086
rect -605 -1126 -547 -1120
rect -413 -1086 -355 -1080
rect -413 -1120 -401 -1086
rect -367 -1120 -355 -1086
rect -413 -1126 -355 -1120
rect -221 -1086 -163 -1080
rect -221 -1120 -209 -1086
rect -175 -1120 -163 -1086
rect -221 -1126 -163 -1120
rect -29 -1086 29 -1080
rect -29 -1120 -17 -1086
rect 17 -1120 29 -1086
rect -29 -1126 29 -1120
rect 163 -1086 221 -1080
rect 163 -1120 175 -1086
rect 209 -1120 221 -1086
rect 163 -1126 221 -1120
rect 355 -1086 413 -1080
rect 355 -1120 367 -1086
rect 401 -1120 413 -1086
rect 355 -1126 413 -1120
rect 547 -1086 605 -1080
rect 547 -1120 559 -1086
rect 593 -1120 605 -1086
rect 547 -1126 605 -1120
rect 739 -1086 797 -1080
rect 739 -1120 751 -1086
rect 785 -1120 797 -1086
rect 739 -1126 797 -1120
rect 931 -1086 989 -1080
rect 931 -1120 943 -1086
rect 977 -1120 989 -1086
rect 931 -1126 989 -1120
<< properties >>
string FIXED_BBOX -1122 -1205 1122 1205
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10.476190476190476 l 0.15 m 1 nf 21 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
