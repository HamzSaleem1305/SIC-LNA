magic
tech sky130A
magscale 1 2
timestamp 1666356932
<< error_p >>
rect -845 1072 -787 1078
rect -653 1072 -595 1078
rect -461 1072 -403 1078
rect -269 1072 -211 1078
rect -77 1072 -19 1078
rect 115 1072 173 1078
rect 307 1072 365 1078
rect 499 1072 557 1078
rect 691 1072 749 1078
rect 883 1072 941 1078
rect -845 1038 -833 1072
rect -653 1038 -641 1072
rect -461 1038 -449 1072
rect -269 1038 -257 1072
rect -77 1038 -65 1072
rect 115 1038 127 1072
rect 307 1038 319 1072
rect 499 1038 511 1072
rect 691 1038 703 1072
rect 883 1038 895 1072
rect -845 1032 -787 1038
rect -653 1032 -595 1038
rect -461 1032 -403 1038
rect -269 1032 -211 1038
rect -77 1032 -19 1038
rect 115 1032 173 1038
rect 307 1032 365 1038
rect 499 1032 557 1038
rect 691 1032 749 1038
rect 883 1032 941 1038
rect -941 -1038 -883 -1032
rect -749 -1038 -691 -1032
rect -557 -1038 -499 -1032
rect -365 -1038 -307 -1032
rect -173 -1038 -115 -1032
rect 19 -1038 77 -1032
rect 211 -1038 269 -1032
rect 403 -1038 461 -1032
rect 595 -1038 653 -1032
rect 787 -1038 845 -1032
rect -941 -1072 -929 -1038
rect -749 -1072 -737 -1038
rect -557 -1072 -545 -1038
rect -365 -1072 -353 -1038
rect -173 -1072 -161 -1038
rect 19 -1072 31 -1038
rect 211 -1072 223 -1038
rect 403 -1072 415 -1038
rect 595 -1072 607 -1038
rect 787 -1072 799 -1038
rect -941 -1078 -883 -1072
rect -749 -1078 -691 -1072
rect -557 -1078 -499 -1072
rect -365 -1078 -307 -1072
rect -173 -1078 -115 -1072
rect 19 -1078 77 -1072
rect 211 -1078 269 -1072
rect 403 -1078 461 -1072
rect 595 -1078 653 -1072
rect 787 -1078 845 -1072
<< pwell >>
rect -1127 -1210 1127 1210
<< nmoslvt >>
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
<< ndiff >>
rect -989 988 -927 1000
rect -989 -988 -977 988
rect -943 -988 -927 988
rect -989 -1000 -927 -988
rect -897 988 -831 1000
rect -897 -988 -881 988
rect -847 -988 -831 988
rect -897 -1000 -831 -988
rect -801 988 -735 1000
rect -801 -988 -785 988
rect -751 -988 -735 988
rect -801 -1000 -735 -988
rect -705 988 -639 1000
rect -705 -988 -689 988
rect -655 -988 -639 988
rect -705 -1000 -639 -988
rect -609 988 -543 1000
rect -609 -988 -593 988
rect -559 -988 -543 988
rect -609 -1000 -543 -988
rect -513 988 -447 1000
rect -513 -988 -497 988
rect -463 -988 -447 988
rect -513 -1000 -447 -988
rect -417 988 -351 1000
rect -417 -988 -401 988
rect -367 -988 -351 988
rect -417 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 417 1000
rect 351 -988 367 988
rect 401 -988 417 988
rect 351 -1000 417 -988
rect 447 988 513 1000
rect 447 -988 463 988
rect 497 -988 513 988
rect 447 -1000 513 -988
rect 543 988 609 1000
rect 543 -988 559 988
rect 593 -988 609 988
rect 543 -1000 609 -988
rect 639 988 705 1000
rect 639 -988 655 988
rect 689 -988 705 988
rect 639 -1000 705 -988
rect 735 988 801 1000
rect 735 -988 751 988
rect 785 -988 801 988
rect 735 -1000 801 -988
rect 831 988 897 1000
rect 831 -988 847 988
rect 881 -988 897 988
rect 831 -1000 897 -988
rect 927 988 989 1000
rect 927 -988 943 988
rect 977 -988 989 988
rect 927 -1000 989 -988
<< ndiffc >>
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
<< psubdiff >>
rect -1091 1140 -995 1174
rect 995 1140 1091 1174
rect -1091 1078 -1057 1140
rect 1057 1078 1091 1140
rect -1091 -1140 -1057 -1078
rect 1057 -1140 1091 -1078
rect -1091 -1174 -995 -1140
rect 995 -1174 1091 -1140
<< psubdiffcont >>
rect -995 1140 995 1174
rect -1091 -1078 -1057 1078
rect 1057 -1078 1091 1078
rect -995 -1174 995 -1140
<< poly >>
rect -849 1072 -783 1088
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -927 1000 -897 1026
rect -849 1022 -783 1038
rect -657 1072 -591 1088
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -831 1000 -801 1022
rect -735 1000 -705 1026
rect -657 1022 -591 1038
rect -465 1072 -399 1088
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -639 1000 -609 1022
rect -543 1000 -513 1026
rect -465 1022 -399 1038
rect -273 1072 -207 1088
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -447 1000 -417 1022
rect -351 1000 -321 1026
rect -273 1022 -207 1038
rect -81 1072 -15 1088
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect -255 1000 -225 1022
rect -159 1000 -129 1026
rect -81 1022 -15 1038
rect 111 1072 177 1088
rect 111 1038 127 1072
rect 161 1038 177 1072
rect -63 1000 -33 1022
rect 33 1000 63 1026
rect 111 1022 177 1038
rect 303 1072 369 1088
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 129 1000 159 1022
rect 225 1000 255 1026
rect 303 1022 369 1038
rect 495 1072 561 1088
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 321 1000 351 1022
rect 417 1000 447 1026
rect 495 1022 561 1038
rect 687 1072 753 1088
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 513 1000 543 1022
rect 609 1000 639 1026
rect 687 1022 753 1038
rect 879 1072 945 1088
rect 879 1038 895 1072
rect 929 1038 945 1072
rect 705 1000 735 1022
rect 801 1000 831 1026
rect 879 1022 945 1038
rect 897 1000 927 1022
rect -927 -1022 -897 -1000
rect -945 -1038 -879 -1022
rect -831 -1026 -801 -1000
rect -735 -1022 -705 -1000
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -945 -1088 -879 -1072
rect -753 -1038 -687 -1022
rect -639 -1026 -609 -1000
rect -543 -1022 -513 -1000
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -753 -1088 -687 -1072
rect -561 -1038 -495 -1022
rect -447 -1026 -417 -1000
rect -351 -1022 -321 -1000
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -561 -1088 -495 -1072
rect -369 -1038 -303 -1022
rect -255 -1026 -225 -1000
rect -159 -1022 -129 -1000
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -369 -1088 -303 -1072
rect -177 -1038 -111 -1022
rect -63 -1026 -33 -1000
rect 33 -1022 63 -1000
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect -177 -1088 -111 -1072
rect 15 -1038 81 -1022
rect 129 -1026 159 -1000
rect 225 -1022 255 -1000
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 15 -1088 81 -1072
rect 207 -1038 273 -1022
rect 321 -1026 351 -1000
rect 417 -1022 447 -1000
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 207 -1088 273 -1072
rect 399 -1038 465 -1022
rect 513 -1026 543 -1000
rect 609 -1022 639 -1000
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 399 -1088 465 -1072
rect 591 -1038 657 -1022
rect 705 -1026 735 -1000
rect 801 -1022 831 -1000
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 591 -1088 657 -1072
rect 783 -1038 849 -1022
rect 897 -1026 927 -1000
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect 783 -1088 849 -1072
<< polycont >>
rect -833 1038 -799 1072
rect -641 1038 -607 1072
rect -449 1038 -415 1072
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect 511 1038 545 1072
rect 703 1038 737 1072
rect 895 1038 929 1072
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
<< locali >>
rect -1091 1140 -995 1174
rect 995 1140 1091 1174
rect -1091 1078 -1057 1140
rect 1057 1078 1091 1140
rect -849 1038 -833 1072
rect -799 1038 -783 1072
rect -657 1038 -641 1072
rect -607 1038 -591 1072
rect -465 1038 -449 1072
rect -415 1038 -399 1072
rect -273 1038 -257 1072
rect -223 1038 -207 1072
rect -81 1038 -65 1072
rect -31 1038 -15 1072
rect 111 1038 127 1072
rect 161 1038 177 1072
rect 303 1038 319 1072
rect 353 1038 369 1072
rect 495 1038 511 1072
rect 545 1038 561 1072
rect 687 1038 703 1072
rect 737 1038 753 1072
rect 879 1038 895 1072
rect 929 1038 945 1072
rect -977 988 -943 1004
rect -977 -1004 -943 -988
rect -881 988 -847 1004
rect -881 -1004 -847 -988
rect -785 988 -751 1004
rect -785 -1004 -751 -988
rect -689 988 -655 1004
rect -689 -1004 -655 -988
rect -593 988 -559 1004
rect -593 -1004 -559 -988
rect -497 988 -463 1004
rect -497 -1004 -463 -988
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect 463 988 497 1004
rect 463 -1004 497 -988
rect 559 988 593 1004
rect 559 -1004 593 -988
rect 655 988 689 1004
rect 655 -1004 689 -988
rect 751 988 785 1004
rect 751 -1004 785 -988
rect 847 988 881 1004
rect 847 -1004 881 -988
rect 943 988 977 1004
rect 943 -1004 977 -988
rect -945 -1072 -929 -1038
rect -895 -1072 -879 -1038
rect -753 -1072 -737 -1038
rect -703 -1072 -687 -1038
rect -561 -1072 -545 -1038
rect -511 -1072 -495 -1038
rect -369 -1072 -353 -1038
rect -319 -1072 -303 -1038
rect -177 -1072 -161 -1038
rect -127 -1072 -111 -1038
rect 15 -1072 31 -1038
rect 65 -1072 81 -1038
rect 207 -1072 223 -1038
rect 257 -1072 273 -1038
rect 399 -1072 415 -1038
rect 449 -1072 465 -1038
rect 591 -1072 607 -1038
rect 641 -1072 657 -1038
rect 783 -1072 799 -1038
rect 833 -1072 849 -1038
rect -1091 -1140 -1057 -1078
rect 1057 -1140 1091 -1078
rect -1091 -1174 -995 -1140
rect 995 -1174 1091 -1140
<< viali >>
rect -833 1038 -799 1072
rect -641 1038 -607 1072
rect -449 1038 -415 1072
rect -257 1038 -223 1072
rect -65 1038 -31 1072
rect 127 1038 161 1072
rect 319 1038 353 1072
rect 511 1038 545 1072
rect 703 1038 737 1072
rect 895 1038 929 1072
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect -929 -1072 -895 -1038
rect -737 -1072 -703 -1038
rect -545 -1072 -511 -1038
rect -353 -1072 -319 -1038
rect -161 -1072 -127 -1038
rect 31 -1072 65 -1038
rect 223 -1072 257 -1038
rect 415 -1072 449 -1038
rect 607 -1072 641 -1038
rect 799 -1072 833 -1038
<< metal1 >>
rect -845 1072 -787 1078
rect -845 1038 -833 1072
rect -799 1038 -787 1072
rect -845 1032 -787 1038
rect -653 1072 -595 1078
rect -653 1038 -641 1072
rect -607 1038 -595 1072
rect -653 1032 -595 1038
rect -461 1072 -403 1078
rect -461 1038 -449 1072
rect -415 1038 -403 1072
rect -461 1032 -403 1038
rect -269 1072 -211 1078
rect -269 1038 -257 1072
rect -223 1038 -211 1072
rect -269 1032 -211 1038
rect -77 1072 -19 1078
rect -77 1038 -65 1072
rect -31 1038 -19 1072
rect -77 1032 -19 1038
rect 115 1072 173 1078
rect 115 1038 127 1072
rect 161 1038 173 1072
rect 115 1032 173 1038
rect 307 1072 365 1078
rect 307 1038 319 1072
rect 353 1038 365 1072
rect 307 1032 365 1038
rect 499 1072 557 1078
rect 499 1038 511 1072
rect 545 1038 557 1072
rect 499 1032 557 1038
rect 691 1072 749 1078
rect 691 1038 703 1072
rect 737 1038 749 1072
rect 691 1032 749 1038
rect 883 1072 941 1078
rect 883 1038 895 1072
rect 929 1038 941 1072
rect 883 1032 941 1038
rect -983 988 -937 1000
rect -983 -988 -977 988
rect -943 -988 -937 988
rect -983 -1000 -937 -988
rect -887 988 -841 1000
rect -887 -988 -881 988
rect -847 -988 -841 988
rect -887 -1000 -841 -988
rect -791 988 -745 1000
rect -791 -988 -785 988
rect -751 -988 -745 988
rect -791 -1000 -745 -988
rect -695 988 -649 1000
rect -695 -988 -689 988
rect -655 -988 -649 988
rect -695 -1000 -649 -988
rect -599 988 -553 1000
rect -599 -988 -593 988
rect -559 -988 -553 988
rect -599 -1000 -553 -988
rect -503 988 -457 1000
rect -503 -988 -497 988
rect -463 -988 -457 988
rect -503 -1000 -457 -988
rect -407 988 -361 1000
rect -407 -988 -401 988
rect -367 -988 -361 988
rect -407 -1000 -361 -988
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect 361 988 407 1000
rect 361 -988 367 988
rect 401 -988 407 988
rect 361 -1000 407 -988
rect 457 988 503 1000
rect 457 -988 463 988
rect 497 -988 503 988
rect 457 -1000 503 -988
rect 553 988 599 1000
rect 553 -988 559 988
rect 593 -988 599 988
rect 553 -1000 599 -988
rect 649 988 695 1000
rect 649 -988 655 988
rect 689 -988 695 988
rect 649 -1000 695 -988
rect 745 988 791 1000
rect 745 -988 751 988
rect 785 -988 791 988
rect 745 -1000 791 -988
rect 841 988 887 1000
rect 841 -988 847 988
rect 881 -988 887 988
rect 841 -1000 887 -988
rect 937 988 983 1000
rect 937 -988 943 988
rect 977 -988 983 988
rect 937 -1000 983 -988
rect -941 -1038 -883 -1032
rect -941 -1072 -929 -1038
rect -895 -1072 -883 -1038
rect -941 -1078 -883 -1072
rect -749 -1038 -691 -1032
rect -749 -1072 -737 -1038
rect -703 -1072 -691 -1038
rect -749 -1078 -691 -1072
rect -557 -1038 -499 -1032
rect -557 -1072 -545 -1038
rect -511 -1072 -499 -1038
rect -557 -1078 -499 -1072
rect -365 -1038 -307 -1032
rect -365 -1072 -353 -1038
rect -319 -1072 -307 -1038
rect -365 -1078 -307 -1072
rect -173 -1038 -115 -1032
rect -173 -1072 -161 -1038
rect -127 -1072 -115 -1038
rect -173 -1078 -115 -1072
rect 19 -1038 77 -1032
rect 19 -1072 31 -1038
rect 65 -1072 77 -1038
rect 19 -1078 77 -1072
rect 211 -1038 269 -1032
rect 211 -1072 223 -1038
rect 257 -1072 269 -1038
rect 211 -1078 269 -1072
rect 403 -1038 461 -1032
rect 403 -1072 415 -1038
rect 449 -1072 461 -1038
rect 403 -1078 461 -1072
rect 595 -1038 653 -1032
rect 595 -1072 607 -1038
rect 641 -1072 653 -1038
rect 595 -1078 653 -1072
rect 787 -1038 845 -1032
rect 787 -1072 799 -1038
rect 833 -1072 845 -1038
rect 787 -1078 845 -1072
<< properties >>
string FIXED_BBOX -1074 -1157 1074 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
