magic
tech sky130A
magscale 1 2
timestamp 1666697857
<< metal5 >>
rect 3550 34719 32561 46719
tri 15550 30719 19550 34719 ne
rect 19550 30719 32561 34719
rect 3550 27343 15550 30719
tri 15550 27343 18926 30719 sw
tri 19550 27343 22926 30719 ne
rect 22926 27343 32561 30719
rect 3550 25319 18926 27343
tri 18926 25319 20950 27343 sw
rect 3550 24119 31550 25319
rect 3550 22095 18926 24119
tri 18926 22095 20950 24119 nw
rect 3550 18719 15550 22095
tri 15550 18719 18926 22095 nw
tri 19550 18719 22926 22095 se
rect 22926 18719 32561 22095
tri 15550 14719 19550 18719 se
rect 19550 14719 32561 18719
rect 3550 2719 32561 14719
<< end >>
