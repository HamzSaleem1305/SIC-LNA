magic
tech sky130A
magscale 1 2
timestamp 1666381508
<< pwell >>
rect -201 -1398 201 1398
<< psubdiff >>
rect -165 1328 -69 1362
rect 69 1328 165 1362
rect -165 1266 -131 1328
rect 131 1266 165 1328
rect -165 -1328 -131 -1266
rect 131 -1328 165 -1266
rect -165 -1362 -69 -1328
rect 69 -1362 165 -1328
<< psubdiffcont >>
rect -69 1328 69 1362
rect -165 -1266 -131 1266
rect 131 -1266 165 1266
rect -69 -1362 69 -1328
<< xpolycontact >>
rect -35 800 35 1232
rect -35 -1232 35 -800
<< ppolyres >>
rect -35 -800 35 800
<< locali >>
rect -165 1328 -69 1362
rect 69 1328 165 1362
rect -165 1266 -131 1328
rect 131 1266 165 1328
rect -165 -1328 -131 -1266
rect 131 -1328 165 -1266
rect -165 -1362 -69 -1328
rect 69 -1362 165 -1328
<< viali >>
rect -19 817 19 1214
rect -19 -1214 19 -817
<< metal1 >>
rect -25 1214 25 1226
rect -25 817 -19 1214
rect 19 817 25 1214
rect -25 805 25 817
rect -25 -817 25 -805
rect -25 -1214 -19 -817
rect 19 -1214 25 -817
rect -25 -1226 25 -1214
<< res0p35 >>
rect -37 -802 37 802
<< properties >>
string FIXED_BBOX -148 -1345 148 1345
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 8.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 7.419k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
