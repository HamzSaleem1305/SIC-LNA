magic
tech sky130A
magscale 1 2
timestamp 1666417074
<< pwell >>
rect -201 -1218 201 1218
<< psubdiff >>
rect -165 1148 -69 1182
rect 69 1148 165 1182
rect -165 1086 -131 1148
rect 131 1086 165 1148
rect -165 -1148 -131 -1086
rect 131 -1148 165 -1086
rect -165 -1182 -69 -1148
rect 69 -1182 165 -1148
<< psubdiffcont >>
rect -69 1148 69 1182
rect -165 -1086 -131 1086
rect 131 -1086 165 1086
rect -69 -1182 69 -1148
<< xpolycontact >>
rect -35 620 35 1052
rect -35 -1052 35 -620
<< ppolyres >>
rect -35 -620 35 620
<< locali >>
rect -165 1148 -69 1182
rect 69 1148 165 1182
rect -165 1086 -131 1148
rect 131 1086 165 1148
rect -165 -1148 -131 -1086
rect 131 -1148 165 -1086
rect -165 -1182 -69 -1148
rect 69 -1182 165 -1148
<< viali >>
rect -19 637 19 1034
rect -19 -1034 19 -637
<< metal1 >>
rect -25 1034 25 1046
rect -25 637 -19 1034
rect 19 637 25 1034
rect -25 625 25 637
rect -25 -637 25 -625
rect -25 -1034 -19 -637
rect 19 -1034 25 -637
rect -25 -1046 25 -1034
<< res0p35 >>
rect -37 -622 37 622
<< properties >>
string FIXED_BBOX -148 -1165 148 1165
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 6.2 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 5.774k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
