** sch_path: /home/shahid/Desktop/EDA/test/lna_extra/xschem4_sic_final/2stage_tb_sym.sch
**.subckt 2stage_tb_sym
C6 Vii net2 10n m=1
VIN4 net1 GND sin 0 3m 2e9 0 0 0
VIN5 Vii net1 sin 0 3m 3e9 0 0 0
VIN2 net3 GND sin 0 3m 2e9 0 0 180
C1 net3 net5 10n m=1
VIN1 net4 GND sin 0 0.005m 2e9 0 0 0
C2 net4 net6 10n m=1
VDD9 0_6 GND 0.6
VDD1 0_75 GND 0.75
VDD2 0_9 GND 0.9
VDD3 1_4 GND 1.4
VDD4 1_5 GND 1.55
VDD5 1_8 GND 1.8
X1 1_8 GND VOUT VOUT1 VOUT2 VTEST1 net2 net5 net6 0_75 1_5 1_4 0_9 0_6 2stage_for_symbol
**** begin user architecture code



.control
tran 1p 20n


print @m.xm15.msky130_fd_pr__nfet_01v8_lvt[id]
print @m.xm14.msky130_fd_pr__nfet_01v8_lvt[id]
print @m.xm16.msky130_fd_pr__pfet_01v8[id]
print @m.xm3.msky130_fd_pr__nfet_01v8_lvt[id]

print @m.xm15.msky130_fd_pr__nfet_01v8_lvt[vth]
print @m.xm14.msky130_fd_pr__nfet_01v8_lvt[vth]
print @m.xm16.msky130_fd_pr__pfet_01v8[vth]
print @m.xm3.msky130_fd_pr__nfet_01v8_lvt[vth]

print @m.xm15.msky130_fd_pr__nfet_01v8_lvt[gm]
print @m.xm14.msky130_fd_pr__nfet_01v8_lvt[gm]
print @m.xm16.msky130_fd_pr__pfet_01v8[gm]
print @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]


#plot v(Vo1nn)
#plot v(Vo1n)
#plot v(VI)
#plot v(Vsi)
#plot v(vo1nn)
spectrum 500MEG 7000MEG 50MEG v(VOUT)
let abc=spectrum 500MEG 7000MEG 50MEG v(VOUT)
plot db(abc)

.endc



.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  2stage_for_symbol.sym # of pins=14
** sym_path: /home/shahid/Desktop/EDA/test/lna_extra/xschem4_sic_final/2stage_for_symbol.sym
** sch_path: /home/shahid/Desktop/EDA/test/lna_extra/xschem4_sic_final/2stage_for_symbol.sch
.subckt 2stage_for_symbol  VDD VSS VOUT VOUT1 VOUT2 VTEST1 VRF VSI1 VSI2 VB0_75 VB1_5 VB1_4 VB0_9
+ VB0_6
*.iopin VRF
*.iopin VSS
*.iopin VB0_75
*.iopin VSI1
*.iopin VDD
*.iopin VOUT1
*.iopin VOUT2
*.iopin VB1_4
*.iopin VB1_5
*.iopin VB0_9
*.iopin VSI2
*.iopin VB0_6
*.iopin VTEST1
*.iopin VOUT
XR4 VB1_5 net1 VSS sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XC5 net1 VOUT1 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XM12 VTEST1 VRF VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=200 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 VTEST1 VRF VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=60 nf=11 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 VOUT1 VB1_4 VTEST1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=80 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net2 net1 VRF VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM16 VRF VB0_75 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 VOUT net5 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=45 nf=9 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 VDD net3 VOUT VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3
XR11 net3 VDD VSS sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XM19 VOUT net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16
XC7 VOUT2 net3 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XR12 VB0_9 net5 VSS sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
XC8 VOUT1 net5 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XR13 VB0_6 net4 VSS sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XR14 net2 VDD VSS sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
XM20 VTEST1 VSI1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=220 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR15 VOUT1 VDD VSS sky130_fd_pr__res_high_po_0p69 L=0.69 mult=8 m=8
XR16 VB0_75 VSI1 VSS sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
XM21 VOUT2 VOUT1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR17 VOUT2 VDD VSS sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
XM22 VOUT VSI2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=80 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR18 VB0_75 VSI2 VSS sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
.ends

.GLOBAL GND
.end
