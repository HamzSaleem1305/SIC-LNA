magic
tech sky130A
magscale 1 2
timestamp 1666377285
<< locali >>
rect 13652 8363 13802 8615
rect 11440 7050 11560 7160
rect 11650 6720 15437 6746
rect 11650 6610 11670 6720
rect 11800 6620 12960 6720
rect 13080 6620 14180 6720
rect 14290 6620 15437 6720
rect 11800 6610 15437 6620
rect 11650 6594 15437 6610
rect 15285 6379 15437 6594
<< viali >>
rect 11670 6610 11800 6720
rect 12960 6620 13080 6720
rect 14180 6620 14290 6720
<< metal1 >>
rect 11650 6720 11830 10020
rect 12480 6980 12660 10020
rect 13382 9000 14670 9073
rect 13382 8870 13455 9000
rect 13380 8810 13460 8870
rect 13790 8810 13870 8870
rect 14597 8695 14670 9000
rect 12480 6860 12500 6980
rect 12630 6860 12660 6980
rect 12480 6840 12660 6860
rect 12715 8382 13389 8495
rect 11650 6610 11670 6720
rect 11800 6610 11830 6720
rect 11650 6590 11830 6610
rect 11860 6678 11956 6683
rect 12715 6678 12828 8382
rect 14131 8143 14318 8518
rect 12985 8119 13099 8137
rect 12985 7892 12998 8119
rect 13081 7892 13099 8119
rect 12985 7880 13099 7892
rect 13448 8121 13531 8137
rect 13448 7892 13459 8121
rect 13519 7892 13531 8121
rect 13448 7882 13531 7892
rect 13850 7888 14318 8143
rect 13850 7887 14278 7888
rect 11860 6670 12828 6678
rect 11860 6575 11872 6670
rect 11936 6575 12828 6670
rect 12940 6720 13100 7290
rect 13448 7229 13609 7330
rect 12940 6620 12960 6720
rect 13080 6620 13100 6720
rect 12940 6600 13100 6620
rect 13360 7185 13470 7190
rect 13360 6770 13474 7185
rect 13788 6978 13877 7191
rect 13788 6852 13800 6978
rect 13859 6852 13877 6978
rect 13788 6840 13877 6852
rect 11860 6565 12828 6575
rect 13360 6570 13370 6770
rect 13460 6570 13474 6770
rect 14160 6720 14320 7270
rect 14593 7170 14949 7427
rect 14160 6620 14180 6720
rect 14290 6620 14320 6720
rect 14160 6594 14320 6620
rect 13360 6560 13474 6570
rect 13367 6559 13474 6560
rect 11851 5725 11946 5738
rect 11851 5606 11864 5725
rect 11933 5606 11946 5725
rect 11851 5593 11946 5606
<< via1 >>
rect 12500 6860 12630 6980
rect 12998 7892 13081 8119
rect 13459 7892 13519 8121
rect 11872 6575 11936 6670
rect 13800 6852 13859 6978
rect 13370 6570 13460 6770
rect 11864 5606 11933 5725
<< metal2 >>
rect 12986 8121 13531 8137
rect 12986 8119 13459 8121
rect 12986 7892 12998 8119
rect 13081 7892 13459 8119
rect 13519 7892 13531 8121
rect 12986 7880 13531 7892
rect 16454 7569 16865 7592
rect 16454 7491 16490 7569
rect 15085 7331 16490 7491
rect 15085 7000 15245 7331
rect 16454 7293 16490 7331
rect 16835 7293 16865 7569
rect 16454 7266 16865 7293
rect 12480 6980 15245 7000
rect 12480 6860 12500 6980
rect 12630 6978 15245 6980
rect 12630 6860 13800 6978
rect 12480 6852 13800 6860
rect 13859 6852 15245 6978
rect 12480 6840 15245 6852
rect 11850 6670 11946 6683
rect 11850 6575 11872 6670
rect 11936 6575 11946 6670
rect 11850 6565 11946 6575
rect 12830 6070 12990 6840
rect 13360 6770 13470 6780
rect 13360 6570 13370 6770
rect 13460 6570 13470 6770
rect 13360 6560 13470 6570
rect 11851 5725 11946 5738
rect 11851 5606 11864 5725
rect 11933 5606 11946 5725
rect 11851 5593 11946 5606
<< via2 >>
rect 16490 7293 16835 7569
rect 11872 6575 11936 6670
rect 13370 6570 13460 6770
rect 11864 5606 11933 5725
<< metal3 >>
rect 16454 7569 16865 7592
rect 16454 7293 16490 7569
rect 16835 7293 16865 7569
rect 16454 7266 16865 7293
rect 16660 6870 16930 6900
rect 16660 6785 16680 6870
rect 13359 6770 16680 6785
rect 11851 6670 11946 6682
rect 11851 6575 11872 6670
rect 11936 6575 11946 6670
rect 11851 5725 11946 6575
rect 13359 6574 13370 6770
rect 13360 6570 13370 6574
rect 13460 6574 16680 6770
rect 13460 6570 13470 6574
rect 13360 6560 13470 6570
rect 16660 6540 16680 6574
rect 16910 6540 16930 6870
rect 16660 6510 16930 6540
rect 11851 5606 11864 5725
rect 11933 5606 11946 5725
rect 11851 5593 11946 5606
<< via3 >>
rect 16490 7293 16835 7569
rect 16680 6540 16910 6870
<< metal4 >>
rect 16454 7569 17572 7591
rect 16454 7293 16490 7569
rect 16835 7293 17572 7569
rect 16454 7266 17572 7293
rect 16660 6871 16930 6900
rect 16660 6538 16676 6871
rect 16916 6538 16930 6871
rect 16660 6510 16930 6538
<< via4 >>
rect 16676 6870 16916 6871
rect 16676 6540 16680 6870
rect 16680 6540 16910 6870
rect 16910 6540 16916 6870
rect 16676 6538 16916 6540
<< metal5 >>
rect 16625 6871 17430 6900
rect 16625 6538 16676 6871
rect 16916 6538 17430 6871
rect 16625 6510 17430 6538
use sky130_fd_pr__cap_mim_m3_2_3HBNLG  XC5
timestamp 1666374491
transform 0 -1 20304 1 0 4217
box -3351 -3101 3373 3101
use sky130_fd_pr__nfet_01v8_lvt_PDNSV3  XM15
timestamp 1666374491
transform 1 0 13421 0 1 8000
box -211 -990 211 990
use sky130_fd_pr__nfet_01v8_lvt_PDNSV3  XM21
timestamp 1666374491
transform 1 0 13831 0 1 8000
box -211 -990 211 990
use sky130_fd_pr__res_high_po_0p35_HCAWEA  XR4
timestamp 1666374491
transform 1 0 14633 0 1 8009
box -201 -998 201 998
use sky130_fd_pr__res_high_po_0p35_SVGS7M  XR14
timestamp 1666374491
transform 1 0 13021 0 1 7658
box -201 -648 201 648
use sky130_fd_pr__res_high_po_0p35_SVGS7M  XR17
timestamp 1666374491
transform 1 0 14241 0 1 7658
box -201 -648 201 648
use sky130_fd_pr__res_high_po_0p69_NCBZCX  sky130_fd_pr__res_high_po_0p69_NCBZCX_0
timestamp 1666374491
transform 0 -1 12157 1 0 8596
box -1586 -667 1586 667
<< labels >>
flabel metal1 14875 7282 14875 7282 0 FreeSans 1600 0 0 0 VB1_5
flabel metal1 14219 8433 14219 8440 0 FreeSans 800 0 0 0 VOUT2
flabel metal3 11889 6510 11889 6510 0 FreeSans 800 0 0 0 VRF
flabel metal2 14941 6915 14941 6915 0 FreeSans 800 0 0 0 VOUT1
flabel locali 12210 6720 12210 6720 0 FreeSans 800 0 0 0 VDD
flabel locali 11470 7100 11470 7100 0 FreeSans 800 0 0 0 VSS
<< end >>
