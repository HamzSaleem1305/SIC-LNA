magic
tech sky130A
timestamp 1640952342
<< error_p >>
rect -54 -525 -25 525
rect 25 -525 54 525
<< nmos >>
rect -25 -525 25 525
<< ndiff >>
rect -54 519 -25 525
rect -54 -519 -48 519
rect -31 -519 -25 519
rect -54 -525 -25 -519
rect 25 519 54 525
rect 25 -519 31 519
rect 48 -519 54 519
rect 25 -525 54 -519
<< ndiffc >>
rect -48 -519 -31 519
rect 31 -519 48 519
<< poly >>
rect -25 525 25 538
rect -25 -538 25 -525
<< locali >>
rect -48 519 -31 527
rect -48 -527 -31 -519
rect 31 519 48 527
rect 31 -527 48 -519
<< viali >>
rect -48 -519 -31 519
rect 31 -519 48 519
<< metal1 >>
rect -51 519 -28 525
rect -51 -519 -48 519
rect -31 -519 -28 519
rect -51 -525 -28 -519
rect 28 519 51 525
rect 28 -519 31 519
rect 48 -519 51 519
rect 28 -525 51 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 10.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
