** sch_path: /home/shahid/Desktop/EDA/test/xschem4_sic_final/CompleteAMP6with50ohms1_ac.sch
**.subckt CompleteAMP6with50ohms1_ac
Vcasc3 net1 GND 1.4
VDD4 net2 GND 1.8
VDD5 net3 GND 1.8
Vbias6 net4 GND 0.75
Vcasc7 net5 GND 1.55
XR1 net5 net6 GND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XC5 net6 Vo1n sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
C6 net8 Vi 10n m=1
XM9 Vo1nn Vi GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=200 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 Vo1nn Vi net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=60 nf=11 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 Vo1n net1 Vo1nn GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=80 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net7 net6 Vi GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 Vi net4 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 Vo2 net13 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=45 nf=9 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net10 net9 Vo2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XR10 net9 net10 GND sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XM16 Vo2 net11 net10 net10 sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16
VDD8 net10 GND 1.8
VDD9 net14 GND 0.6
XC7 Vo1p net9 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
Vcasc10 net12 GND 0.9
XR11 net12 net13 GND sky130_fd_pr__res_high_po_0p35 L=8 mult=1 m=1
XC8 Vo1n net13 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XR12 net14 net11 GND sky130_fd_pr__res_high_po_0p35 L=15 mult=1 m=1
XR14 net7 net2 GND sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
XM1 Vo1nn GND GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=220 nf=20 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VIN3 net15 GND 0.75
VIN4 Vii GND 0 ac 1m
XR13 Vo1n net2 GND sky130_fd_pr__res_high_po_0p69 L=0.69 mult=8 m=8
XR2 net15 GND GND sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
XM2 Vo1p Vo1n GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR3 Vo1p net2 GND sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
R4 Vii net8 50 m=1
XM22 Vo2 GND GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=80 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net10 net16 Vo2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=100 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR5 net16 net10 GND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XC1 Vo2 net16 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XR6 GND Vo2 GND sky130_fd_pr__res_high_po_0p35 L=0.5 mult=1 m=1
**** begin user architecture code

.lib /home/shahid/OSPDKs/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.control
ac dec 100 0.1G 10G
plot db(v(vo2)/v(vii))
let Zo=50;
let Zin=v(vi)/-i(VIN4)
Let S11=mag( (Zin-Zo)/(Zin+Zo) )
plot db(S11)
WRDATA S11.csv db(S11)
plot mag(Zin);

set sqrnoise
noise v(Vo2) VIN4 dec 40 1G 10G
setplot noise1
let Fn=inoise_spectrum/(8.3e-19)
let NFn=db(Fn) / 2
plot NFn


.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
