magic
tech sky130B
magscale 1 2
timestamp 1667060080
<< nwell >>
rect 15680 20970 16302 23408
rect 16942 13724 17564 16162
<< pwell >>
rect 12890 24686 17066 24772
rect 12890 24476 12976 24686
rect 16980 24476 17066 24686
rect 12890 24390 17066 24476
rect 16522 24240 17066 24390
rect 12920 24006 14896 24092
rect 12920 23796 13006 24006
rect 14810 23796 14896 24006
rect 12920 23710 14896 23796
rect 13830 22226 14912 23350
rect 13330 22140 14912 22226
rect 13330 21036 13416 22140
rect 13626 21036 14912 22140
rect 13330 20950 14912 21036
rect 15150 23300 15532 23386
rect 15150 21056 15236 23300
rect 15446 21056 15532 23300
rect 15150 20970 15532 21056
rect 16522 21840 17796 24240
rect 16630 21420 17012 21506
rect 13156 19800 14470 19886
rect 13156 16820 13242 19800
rect 14384 18010 14470 19800
rect 14690 18960 15676 20646
rect 15850 18960 16452 20160
rect 16630 18816 16716 21420
rect 16926 18816 17012 21420
rect 16630 18730 17012 18816
rect 17240 21440 17622 21526
rect 14876 18010 15688 18694
rect 16098 18625 16480 18711
rect 16098 18010 16184 18625
rect 14384 17924 16184 18010
rect 14384 16820 14572 17924
rect 14782 16820 15792 17924
rect 16002 16821 16184 17924
rect 16394 16821 16480 18625
rect 16660 18140 17006 18486
rect 17240 17436 17326 21440
rect 17536 17436 17622 21440
rect 17240 17350 17622 17436
rect 16002 16820 16480 16821
rect 13156 16735 16480 16820
rect 13156 16734 16088 16735
rect 13432 13616 13834 15664
rect 14282 13616 15364 16104
rect 15992 16034 16374 16120
rect 15992 13790 16078 16034
rect 16288 13790 16374 16034
rect 15992 13616 16374 13790
rect 13048 13429 17896 13616
rect 13048 13096 13235 13429
rect 17702 13096 17896 13429
rect 13048 11044 17896 13096
rect 13048 10764 13235 11044
rect 17702 10764 17896 11044
rect 13048 10584 17896 10764
<< pmos >>
rect 15880 21189 15910 23189
rect 15976 21189 16006 23189
rect 16072 21189 16102 23189
rect 17142 13943 17172 15943
rect 17238 13943 17268 15943
rect 17334 13943 17364 15943
<< nmoslvt >>
rect 14020 21150 14050 23150
rect 14116 21150 14146 23150
rect 14212 21150 14242 23150
rect 14308 21150 14338 23150
rect 14404 21150 14434 23150
rect 14500 21150 14530 23150
rect 14596 21150 14626 23150
rect 14692 21150 14722 23150
rect 16712 22040 16742 24040
rect 16808 22040 16838 24040
rect 16904 22040 16934 24040
rect 17000 22040 17030 24040
rect 17096 22040 17126 24040
rect 17192 22040 17222 24040
rect 17288 22040 17318 24040
rect 17384 22040 17414 24040
rect 17480 22040 17510 24040
rect 17576 22040 17606 24040
rect 14880 19160 14910 20446
rect 14976 19160 15006 20446
rect 15072 19160 15102 20446
rect 15168 19160 15198 20446
rect 15264 19160 15294 20446
rect 15360 19160 15390 20446
rect 15456 19160 15486 20446
rect 16040 19160 16070 19960
rect 16136 19160 16166 19960
rect 16232 19160 16262 19960
rect 15062 16934 15092 18494
rect 15472 16934 15502 18494
rect 13618 13904 13648 15464
rect 14472 13904 14502 15904
rect 14568 13904 14598 15904
rect 14664 13904 14694 15904
rect 14760 13904 14790 15904
rect 14856 13904 14886 15904
rect 14952 13904 14982 15904
rect 15048 13904 15078 15904
rect 15144 13904 15174 15904
rect 13480 11070 13510 13070
rect 13568 11070 13598 13070
rect 13656 11070 13686 13070
rect 13744 11070 13774 13070
rect 13832 11070 13862 13070
rect 13920 11070 13950 13070
rect 14008 11070 14038 13070
rect 14096 11070 14126 13070
rect 14184 11070 14214 13070
rect 14272 11070 14302 13070
rect 14360 11070 14390 13070
rect 14448 11070 14478 13070
rect 14536 11070 14566 13070
rect 14624 11070 14654 13070
rect 14712 11070 14742 13070
rect 14800 11070 14830 13070
rect 14888 11070 14918 13070
rect 14976 11070 15006 13070
rect 15064 11070 15094 13070
rect 15152 11070 15182 13070
rect 15240 11070 15270 13070
rect 15328 11070 15358 13070
rect 15416 11070 15446 13070
rect 15504 11070 15534 13070
rect 15592 11070 15622 13070
rect 15680 11070 15710 13070
rect 15768 11070 15798 13070
rect 15856 11070 15886 13070
rect 15944 11070 15974 13070
rect 16032 11070 16062 13070
rect 16120 11070 16150 13070
rect 16208 11070 16238 13070
rect 16296 11070 16326 13070
rect 16384 11070 16414 13070
rect 16472 11070 16502 13070
rect 16560 11070 16590 13070
rect 16648 11070 16678 13070
rect 16736 11070 16766 13070
rect 16824 11070 16854 13070
rect 16912 11070 16942 13070
rect 17000 11070 17030 13070
rect 17088 11070 17118 13070
rect 17176 11070 17206 13070
rect 17264 11070 17294 13070
rect 17352 11070 17382 13070
rect 17440 11070 17470 13070
<< ndiff >>
rect 13958 23119 14020 23150
rect 13958 23085 13970 23119
rect 14004 23085 14020 23119
rect 13958 23051 14020 23085
rect 13958 23017 13970 23051
rect 14004 23017 14020 23051
rect 13958 22983 14020 23017
rect 13958 22949 13970 22983
rect 14004 22949 14020 22983
rect 13958 22915 14020 22949
rect 13958 22881 13970 22915
rect 14004 22881 14020 22915
rect 13958 22847 14020 22881
rect 13958 22813 13970 22847
rect 14004 22813 14020 22847
rect 13958 22779 14020 22813
rect 13958 22745 13970 22779
rect 14004 22745 14020 22779
rect 13958 22711 14020 22745
rect 13958 22677 13970 22711
rect 14004 22677 14020 22711
rect 13958 22643 14020 22677
rect 13958 22609 13970 22643
rect 14004 22609 14020 22643
rect 13958 22575 14020 22609
rect 13958 22541 13970 22575
rect 14004 22541 14020 22575
rect 13958 22507 14020 22541
rect 13958 22473 13970 22507
rect 14004 22473 14020 22507
rect 13958 22439 14020 22473
rect 13958 22405 13970 22439
rect 14004 22405 14020 22439
rect 13958 22371 14020 22405
rect 13958 22337 13970 22371
rect 14004 22337 14020 22371
rect 13958 22303 14020 22337
rect 13958 22269 13970 22303
rect 14004 22269 14020 22303
rect 13958 22235 14020 22269
rect 13958 22201 13970 22235
rect 14004 22201 14020 22235
rect 13958 22167 14020 22201
rect 13958 22133 13970 22167
rect 14004 22133 14020 22167
rect 13958 22099 14020 22133
rect 13958 22065 13970 22099
rect 14004 22065 14020 22099
rect 13958 22031 14020 22065
rect 13958 21997 13970 22031
rect 14004 21997 14020 22031
rect 13958 21963 14020 21997
rect 13958 21929 13970 21963
rect 14004 21929 14020 21963
rect 13958 21895 14020 21929
rect 13958 21861 13970 21895
rect 14004 21861 14020 21895
rect 13958 21827 14020 21861
rect 13958 21793 13970 21827
rect 14004 21793 14020 21827
rect 13958 21759 14020 21793
rect 13958 21725 13970 21759
rect 14004 21725 14020 21759
rect 13958 21691 14020 21725
rect 13958 21657 13970 21691
rect 14004 21657 14020 21691
rect 13958 21623 14020 21657
rect 13958 21589 13970 21623
rect 14004 21589 14020 21623
rect 13958 21555 14020 21589
rect 13958 21521 13970 21555
rect 14004 21521 14020 21555
rect 13958 21487 14020 21521
rect 13958 21453 13970 21487
rect 14004 21453 14020 21487
rect 13958 21419 14020 21453
rect 13958 21385 13970 21419
rect 14004 21385 14020 21419
rect 13958 21351 14020 21385
rect 13958 21317 13970 21351
rect 14004 21317 14020 21351
rect 13958 21283 14020 21317
rect 13958 21249 13970 21283
rect 14004 21249 14020 21283
rect 13958 21215 14020 21249
rect 13958 21181 13970 21215
rect 14004 21181 14020 21215
rect 13958 21150 14020 21181
rect 14050 23119 14116 23150
rect 14050 23085 14066 23119
rect 14100 23085 14116 23119
rect 14050 23051 14116 23085
rect 14050 23017 14066 23051
rect 14100 23017 14116 23051
rect 14050 22983 14116 23017
rect 14050 22949 14066 22983
rect 14100 22949 14116 22983
rect 14050 22915 14116 22949
rect 14050 22881 14066 22915
rect 14100 22881 14116 22915
rect 14050 22847 14116 22881
rect 14050 22813 14066 22847
rect 14100 22813 14116 22847
rect 14050 22779 14116 22813
rect 14050 22745 14066 22779
rect 14100 22745 14116 22779
rect 14050 22711 14116 22745
rect 14050 22677 14066 22711
rect 14100 22677 14116 22711
rect 14050 22643 14116 22677
rect 14050 22609 14066 22643
rect 14100 22609 14116 22643
rect 14050 22575 14116 22609
rect 14050 22541 14066 22575
rect 14100 22541 14116 22575
rect 14050 22507 14116 22541
rect 14050 22473 14066 22507
rect 14100 22473 14116 22507
rect 14050 22439 14116 22473
rect 14050 22405 14066 22439
rect 14100 22405 14116 22439
rect 14050 22371 14116 22405
rect 14050 22337 14066 22371
rect 14100 22337 14116 22371
rect 14050 22303 14116 22337
rect 14050 22269 14066 22303
rect 14100 22269 14116 22303
rect 14050 22235 14116 22269
rect 14050 22201 14066 22235
rect 14100 22201 14116 22235
rect 14050 22167 14116 22201
rect 14050 22133 14066 22167
rect 14100 22133 14116 22167
rect 14050 22099 14116 22133
rect 14050 22065 14066 22099
rect 14100 22065 14116 22099
rect 14050 22031 14116 22065
rect 14050 21997 14066 22031
rect 14100 21997 14116 22031
rect 14050 21963 14116 21997
rect 14050 21929 14066 21963
rect 14100 21929 14116 21963
rect 14050 21895 14116 21929
rect 14050 21861 14066 21895
rect 14100 21861 14116 21895
rect 14050 21827 14116 21861
rect 14050 21793 14066 21827
rect 14100 21793 14116 21827
rect 14050 21759 14116 21793
rect 14050 21725 14066 21759
rect 14100 21725 14116 21759
rect 14050 21691 14116 21725
rect 14050 21657 14066 21691
rect 14100 21657 14116 21691
rect 14050 21623 14116 21657
rect 14050 21589 14066 21623
rect 14100 21589 14116 21623
rect 14050 21555 14116 21589
rect 14050 21521 14066 21555
rect 14100 21521 14116 21555
rect 14050 21487 14116 21521
rect 14050 21453 14066 21487
rect 14100 21453 14116 21487
rect 14050 21419 14116 21453
rect 14050 21385 14066 21419
rect 14100 21385 14116 21419
rect 14050 21351 14116 21385
rect 14050 21317 14066 21351
rect 14100 21317 14116 21351
rect 14050 21283 14116 21317
rect 14050 21249 14066 21283
rect 14100 21249 14116 21283
rect 14050 21215 14116 21249
rect 14050 21181 14066 21215
rect 14100 21181 14116 21215
rect 14050 21150 14116 21181
rect 14146 23119 14212 23150
rect 14146 23085 14162 23119
rect 14196 23085 14212 23119
rect 14146 23051 14212 23085
rect 14146 23017 14162 23051
rect 14196 23017 14212 23051
rect 14146 22983 14212 23017
rect 14146 22949 14162 22983
rect 14196 22949 14212 22983
rect 14146 22915 14212 22949
rect 14146 22881 14162 22915
rect 14196 22881 14212 22915
rect 14146 22847 14212 22881
rect 14146 22813 14162 22847
rect 14196 22813 14212 22847
rect 14146 22779 14212 22813
rect 14146 22745 14162 22779
rect 14196 22745 14212 22779
rect 14146 22711 14212 22745
rect 14146 22677 14162 22711
rect 14196 22677 14212 22711
rect 14146 22643 14212 22677
rect 14146 22609 14162 22643
rect 14196 22609 14212 22643
rect 14146 22575 14212 22609
rect 14146 22541 14162 22575
rect 14196 22541 14212 22575
rect 14146 22507 14212 22541
rect 14146 22473 14162 22507
rect 14196 22473 14212 22507
rect 14146 22439 14212 22473
rect 14146 22405 14162 22439
rect 14196 22405 14212 22439
rect 14146 22371 14212 22405
rect 14146 22337 14162 22371
rect 14196 22337 14212 22371
rect 14146 22303 14212 22337
rect 14146 22269 14162 22303
rect 14196 22269 14212 22303
rect 14146 22235 14212 22269
rect 14146 22201 14162 22235
rect 14196 22201 14212 22235
rect 14146 22167 14212 22201
rect 14146 22133 14162 22167
rect 14196 22133 14212 22167
rect 14146 22099 14212 22133
rect 14146 22065 14162 22099
rect 14196 22065 14212 22099
rect 14146 22031 14212 22065
rect 14146 21997 14162 22031
rect 14196 21997 14212 22031
rect 14146 21963 14212 21997
rect 14146 21929 14162 21963
rect 14196 21929 14212 21963
rect 14146 21895 14212 21929
rect 14146 21861 14162 21895
rect 14196 21861 14212 21895
rect 14146 21827 14212 21861
rect 14146 21793 14162 21827
rect 14196 21793 14212 21827
rect 14146 21759 14212 21793
rect 14146 21725 14162 21759
rect 14196 21725 14212 21759
rect 14146 21691 14212 21725
rect 14146 21657 14162 21691
rect 14196 21657 14212 21691
rect 14146 21623 14212 21657
rect 14146 21589 14162 21623
rect 14196 21589 14212 21623
rect 14146 21555 14212 21589
rect 14146 21521 14162 21555
rect 14196 21521 14212 21555
rect 14146 21487 14212 21521
rect 14146 21453 14162 21487
rect 14196 21453 14212 21487
rect 14146 21419 14212 21453
rect 14146 21385 14162 21419
rect 14196 21385 14212 21419
rect 14146 21351 14212 21385
rect 14146 21317 14162 21351
rect 14196 21317 14212 21351
rect 14146 21283 14212 21317
rect 14146 21249 14162 21283
rect 14196 21249 14212 21283
rect 14146 21215 14212 21249
rect 14146 21181 14162 21215
rect 14196 21181 14212 21215
rect 14146 21150 14212 21181
rect 14242 23119 14308 23150
rect 14242 23085 14258 23119
rect 14292 23085 14308 23119
rect 14242 23051 14308 23085
rect 14242 23017 14258 23051
rect 14292 23017 14308 23051
rect 14242 22983 14308 23017
rect 14242 22949 14258 22983
rect 14292 22949 14308 22983
rect 14242 22915 14308 22949
rect 14242 22881 14258 22915
rect 14292 22881 14308 22915
rect 14242 22847 14308 22881
rect 14242 22813 14258 22847
rect 14292 22813 14308 22847
rect 14242 22779 14308 22813
rect 14242 22745 14258 22779
rect 14292 22745 14308 22779
rect 14242 22711 14308 22745
rect 14242 22677 14258 22711
rect 14292 22677 14308 22711
rect 14242 22643 14308 22677
rect 14242 22609 14258 22643
rect 14292 22609 14308 22643
rect 14242 22575 14308 22609
rect 14242 22541 14258 22575
rect 14292 22541 14308 22575
rect 14242 22507 14308 22541
rect 14242 22473 14258 22507
rect 14292 22473 14308 22507
rect 14242 22439 14308 22473
rect 14242 22405 14258 22439
rect 14292 22405 14308 22439
rect 14242 22371 14308 22405
rect 14242 22337 14258 22371
rect 14292 22337 14308 22371
rect 14242 22303 14308 22337
rect 14242 22269 14258 22303
rect 14292 22269 14308 22303
rect 14242 22235 14308 22269
rect 14242 22201 14258 22235
rect 14292 22201 14308 22235
rect 14242 22167 14308 22201
rect 14242 22133 14258 22167
rect 14292 22133 14308 22167
rect 14242 22099 14308 22133
rect 14242 22065 14258 22099
rect 14292 22065 14308 22099
rect 14242 22031 14308 22065
rect 14242 21997 14258 22031
rect 14292 21997 14308 22031
rect 14242 21963 14308 21997
rect 14242 21929 14258 21963
rect 14292 21929 14308 21963
rect 14242 21895 14308 21929
rect 14242 21861 14258 21895
rect 14292 21861 14308 21895
rect 14242 21827 14308 21861
rect 14242 21793 14258 21827
rect 14292 21793 14308 21827
rect 14242 21759 14308 21793
rect 14242 21725 14258 21759
rect 14292 21725 14308 21759
rect 14242 21691 14308 21725
rect 14242 21657 14258 21691
rect 14292 21657 14308 21691
rect 14242 21623 14308 21657
rect 14242 21589 14258 21623
rect 14292 21589 14308 21623
rect 14242 21555 14308 21589
rect 14242 21521 14258 21555
rect 14292 21521 14308 21555
rect 14242 21487 14308 21521
rect 14242 21453 14258 21487
rect 14292 21453 14308 21487
rect 14242 21419 14308 21453
rect 14242 21385 14258 21419
rect 14292 21385 14308 21419
rect 14242 21351 14308 21385
rect 14242 21317 14258 21351
rect 14292 21317 14308 21351
rect 14242 21283 14308 21317
rect 14242 21249 14258 21283
rect 14292 21249 14308 21283
rect 14242 21215 14308 21249
rect 14242 21181 14258 21215
rect 14292 21181 14308 21215
rect 14242 21150 14308 21181
rect 14338 23119 14404 23150
rect 14338 23085 14354 23119
rect 14388 23085 14404 23119
rect 14338 23051 14404 23085
rect 14338 23017 14354 23051
rect 14388 23017 14404 23051
rect 14338 22983 14404 23017
rect 14338 22949 14354 22983
rect 14388 22949 14404 22983
rect 14338 22915 14404 22949
rect 14338 22881 14354 22915
rect 14388 22881 14404 22915
rect 14338 22847 14404 22881
rect 14338 22813 14354 22847
rect 14388 22813 14404 22847
rect 14338 22779 14404 22813
rect 14338 22745 14354 22779
rect 14388 22745 14404 22779
rect 14338 22711 14404 22745
rect 14338 22677 14354 22711
rect 14388 22677 14404 22711
rect 14338 22643 14404 22677
rect 14338 22609 14354 22643
rect 14388 22609 14404 22643
rect 14338 22575 14404 22609
rect 14338 22541 14354 22575
rect 14388 22541 14404 22575
rect 14338 22507 14404 22541
rect 14338 22473 14354 22507
rect 14388 22473 14404 22507
rect 14338 22439 14404 22473
rect 14338 22405 14354 22439
rect 14388 22405 14404 22439
rect 14338 22371 14404 22405
rect 14338 22337 14354 22371
rect 14388 22337 14404 22371
rect 14338 22303 14404 22337
rect 14338 22269 14354 22303
rect 14388 22269 14404 22303
rect 14338 22235 14404 22269
rect 14338 22201 14354 22235
rect 14388 22201 14404 22235
rect 14338 22167 14404 22201
rect 14338 22133 14354 22167
rect 14388 22133 14404 22167
rect 14338 22099 14404 22133
rect 14338 22065 14354 22099
rect 14388 22065 14404 22099
rect 14338 22031 14404 22065
rect 14338 21997 14354 22031
rect 14388 21997 14404 22031
rect 14338 21963 14404 21997
rect 14338 21929 14354 21963
rect 14388 21929 14404 21963
rect 14338 21895 14404 21929
rect 14338 21861 14354 21895
rect 14388 21861 14404 21895
rect 14338 21827 14404 21861
rect 14338 21793 14354 21827
rect 14388 21793 14404 21827
rect 14338 21759 14404 21793
rect 14338 21725 14354 21759
rect 14388 21725 14404 21759
rect 14338 21691 14404 21725
rect 14338 21657 14354 21691
rect 14388 21657 14404 21691
rect 14338 21623 14404 21657
rect 14338 21589 14354 21623
rect 14388 21589 14404 21623
rect 14338 21555 14404 21589
rect 14338 21521 14354 21555
rect 14388 21521 14404 21555
rect 14338 21487 14404 21521
rect 14338 21453 14354 21487
rect 14388 21453 14404 21487
rect 14338 21419 14404 21453
rect 14338 21385 14354 21419
rect 14388 21385 14404 21419
rect 14338 21351 14404 21385
rect 14338 21317 14354 21351
rect 14388 21317 14404 21351
rect 14338 21283 14404 21317
rect 14338 21249 14354 21283
rect 14388 21249 14404 21283
rect 14338 21215 14404 21249
rect 14338 21181 14354 21215
rect 14388 21181 14404 21215
rect 14338 21150 14404 21181
rect 14434 23119 14500 23150
rect 14434 23085 14450 23119
rect 14484 23085 14500 23119
rect 14434 23051 14500 23085
rect 14434 23017 14450 23051
rect 14484 23017 14500 23051
rect 14434 22983 14500 23017
rect 14434 22949 14450 22983
rect 14484 22949 14500 22983
rect 14434 22915 14500 22949
rect 14434 22881 14450 22915
rect 14484 22881 14500 22915
rect 14434 22847 14500 22881
rect 14434 22813 14450 22847
rect 14484 22813 14500 22847
rect 14434 22779 14500 22813
rect 14434 22745 14450 22779
rect 14484 22745 14500 22779
rect 14434 22711 14500 22745
rect 14434 22677 14450 22711
rect 14484 22677 14500 22711
rect 14434 22643 14500 22677
rect 14434 22609 14450 22643
rect 14484 22609 14500 22643
rect 14434 22575 14500 22609
rect 14434 22541 14450 22575
rect 14484 22541 14500 22575
rect 14434 22507 14500 22541
rect 14434 22473 14450 22507
rect 14484 22473 14500 22507
rect 14434 22439 14500 22473
rect 14434 22405 14450 22439
rect 14484 22405 14500 22439
rect 14434 22371 14500 22405
rect 14434 22337 14450 22371
rect 14484 22337 14500 22371
rect 14434 22303 14500 22337
rect 14434 22269 14450 22303
rect 14484 22269 14500 22303
rect 14434 22235 14500 22269
rect 14434 22201 14450 22235
rect 14484 22201 14500 22235
rect 14434 22167 14500 22201
rect 14434 22133 14450 22167
rect 14484 22133 14500 22167
rect 14434 22099 14500 22133
rect 14434 22065 14450 22099
rect 14484 22065 14500 22099
rect 14434 22031 14500 22065
rect 14434 21997 14450 22031
rect 14484 21997 14500 22031
rect 14434 21963 14500 21997
rect 14434 21929 14450 21963
rect 14484 21929 14500 21963
rect 14434 21895 14500 21929
rect 14434 21861 14450 21895
rect 14484 21861 14500 21895
rect 14434 21827 14500 21861
rect 14434 21793 14450 21827
rect 14484 21793 14500 21827
rect 14434 21759 14500 21793
rect 14434 21725 14450 21759
rect 14484 21725 14500 21759
rect 14434 21691 14500 21725
rect 14434 21657 14450 21691
rect 14484 21657 14500 21691
rect 14434 21623 14500 21657
rect 14434 21589 14450 21623
rect 14484 21589 14500 21623
rect 14434 21555 14500 21589
rect 14434 21521 14450 21555
rect 14484 21521 14500 21555
rect 14434 21487 14500 21521
rect 14434 21453 14450 21487
rect 14484 21453 14500 21487
rect 14434 21419 14500 21453
rect 14434 21385 14450 21419
rect 14484 21385 14500 21419
rect 14434 21351 14500 21385
rect 14434 21317 14450 21351
rect 14484 21317 14500 21351
rect 14434 21283 14500 21317
rect 14434 21249 14450 21283
rect 14484 21249 14500 21283
rect 14434 21215 14500 21249
rect 14434 21181 14450 21215
rect 14484 21181 14500 21215
rect 14434 21150 14500 21181
rect 14530 23119 14596 23150
rect 14530 23085 14546 23119
rect 14580 23085 14596 23119
rect 14530 23051 14596 23085
rect 14530 23017 14546 23051
rect 14580 23017 14596 23051
rect 14530 22983 14596 23017
rect 14530 22949 14546 22983
rect 14580 22949 14596 22983
rect 14530 22915 14596 22949
rect 14530 22881 14546 22915
rect 14580 22881 14596 22915
rect 14530 22847 14596 22881
rect 14530 22813 14546 22847
rect 14580 22813 14596 22847
rect 14530 22779 14596 22813
rect 14530 22745 14546 22779
rect 14580 22745 14596 22779
rect 14530 22711 14596 22745
rect 14530 22677 14546 22711
rect 14580 22677 14596 22711
rect 14530 22643 14596 22677
rect 14530 22609 14546 22643
rect 14580 22609 14596 22643
rect 14530 22575 14596 22609
rect 14530 22541 14546 22575
rect 14580 22541 14596 22575
rect 14530 22507 14596 22541
rect 14530 22473 14546 22507
rect 14580 22473 14596 22507
rect 14530 22439 14596 22473
rect 14530 22405 14546 22439
rect 14580 22405 14596 22439
rect 14530 22371 14596 22405
rect 14530 22337 14546 22371
rect 14580 22337 14596 22371
rect 14530 22303 14596 22337
rect 14530 22269 14546 22303
rect 14580 22269 14596 22303
rect 14530 22235 14596 22269
rect 14530 22201 14546 22235
rect 14580 22201 14596 22235
rect 14530 22167 14596 22201
rect 14530 22133 14546 22167
rect 14580 22133 14596 22167
rect 14530 22099 14596 22133
rect 14530 22065 14546 22099
rect 14580 22065 14596 22099
rect 14530 22031 14596 22065
rect 14530 21997 14546 22031
rect 14580 21997 14596 22031
rect 14530 21963 14596 21997
rect 14530 21929 14546 21963
rect 14580 21929 14596 21963
rect 14530 21895 14596 21929
rect 14530 21861 14546 21895
rect 14580 21861 14596 21895
rect 14530 21827 14596 21861
rect 14530 21793 14546 21827
rect 14580 21793 14596 21827
rect 14530 21759 14596 21793
rect 14530 21725 14546 21759
rect 14580 21725 14596 21759
rect 14530 21691 14596 21725
rect 14530 21657 14546 21691
rect 14580 21657 14596 21691
rect 14530 21623 14596 21657
rect 14530 21589 14546 21623
rect 14580 21589 14596 21623
rect 14530 21555 14596 21589
rect 14530 21521 14546 21555
rect 14580 21521 14596 21555
rect 14530 21487 14596 21521
rect 14530 21453 14546 21487
rect 14580 21453 14596 21487
rect 14530 21419 14596 21453
rect 14530 21385 14546 21419
rect 14580 21385 14596 21419
rect 14530 21351 14596 21385
rect 14530 21317 14546 21351
rect 14580 21317 14596 21351
rect 14530 21283 14596 21317
rect 14530 21249 14546 21283
rect 14580 21249 14596 21283
rect 14530 21215 14596 21249
rect 14530 21181 14546 21215
rect 14580 21181 14596 21215
rect 14530 21150 14596 21181
rect 14626 23119 14692 23150
rect 14626 23085 14642 23119
rect 14676 23085 14692 23119
rect 14626 23051 14692 23085
rect 14626 23017 14642 23051
rect 14676 23017 14692 23051
rect 14626 22983 14692 23017
rect 14626 22949 14642 22983
rect 14676 22949 14692 22983
rect 14626 22915 14692 22949
rect 14626 22881 14642 22915
rect 14676 22881 14692 22915
rect 14626 22847 14692 22881
rect 14626 22813 14642 22847
rect 14676 22813 14692 22847
rect 14626 22779 14692 22813
rect 14626 22745 14642 22779
rect 14676 22745 14692 22779
rect 14626 22711 14692 22745
rect 14626 22677 14642 22711
rect 14676 22677 14692 22711
rect 14626 22643 14692 22677
rect 14626 22609 14642 22643
rect 14676 22609 14692 22643
rect 14626 22575 14692 22609
rect 14626 22541 14642 22575
rect 14676 22541 14692 22575
rect 14626 22507 14692 22541
rect 14626 22473 14642 22507
rect 14676 22473 14692 22507
rect 14626 22439 14692 22473
rect 14626 22405 14642 22439
rect 14676 22405 14692 22439
rect 14626 22371 14692 22405
rect 14626 22337 14642 22371
rect 14676 22337 14692 22371
rect 14626 22303 14692 22337
rect 14626 22269 14642 22303
rect 14676 22269 14692 22303
rect 14626 22235 14692 22269
rect 14626 22201 14642 22235
rect 14676 22201 14692 22235
rect 14626 22167 14692 22201
rect 14626 22133 14642 22167
rect 14676 22133 14692 22167
rect 14626 22099 14692 22133
rect 14626 22065 14642 22099
rect 14676 22065 14692 22099
rect 14626 22031 14692 22065
rect 14626 21997 14642 22031
rect 14676 21997 14692 22031
rect 14626 21963 14692 21997
rect 14626 21929 14642 21963
rect 14676 21929 14692 21963
rect 14626 21895 14692 21929
rect 14626 21861 14642 21895
rect 14676 21861 14692 21895
rect 14626 21827 14692 21861
rect 14626 21793 14642 21827
rect 14676 21793 14692 21827
rect 14626 21759 14692 21793
rect 14626 21725 14642 21759
rect 14676 21725 14692 21759
rect 14626 21691 14692 21725
rect 14626 21657 14642 21691
rect 14676 21657 14692 21691
rect 14626 21623 14692 21657
rect 14626 21589 14642 21623
rect 14676 21589 14692 21623
rect 14626 21555 14692 21589
rect 14626 21521 14642 21555
rect 14676 21521 14692 21555
rect 14626 21487 14692 21521
rect 14626 21453 14642 21487
rect 14676 21453 14692 21487
rect 14626 21419 14692 21453
rect 14626 21385 14642 21419
rect 14676 21385 14692 21419
rect 14626 21351 14692 21385
rect 14626 21317 14642 21351
rect 14676 21317 14692 21351
rect 14626 21283 14692 21317
rect 14626 21249 14642 21283
rect 14676 21249 14692 21283
rect 14626 21215 14692 21249
rect 14626 21181 14642 21215
rect 14676 21181 14692 21215
rect 14626 21150 14692 21181
rect 14722 23119 14784 23150
rect 14722 23085 14738 23119
rect 14772 23085 14784 23119
rect 14722 23051 14784 23085
rect 14722 23017 14738 23051
rect 14772 23017 14784 23051
rect 14722 22983 14784 23017
rect 14722 22949 14738 22983
rect 14772 22949 14784 22983
rect 14722 22915 14784 22949
rect 14722 22881 14738 22915
rect 14772 22881 14784 22915
rect 14722 22847 14784 22881
rect 14722 22813 14738 22847
rect 14772 22813 14784 22847
rect 14722 22779 14784 22813
rect 14722 22745 14738 22779
rect 14772 22745 14784 22779
rect 14722 22711 14784 22745
rect 14722 22677 14738 22711
rect 14772 22677 14784 22711
rect 14722 22643 14784 22677
rect 14722 22609 14738 22643
rect 14772 22609 14784 22643
rect 14722 22575 14784 22609
rect 14722 22541 14738 22575
rect 14772 22541 14784 22575
rect 14722 22507 14784 22541
rect 14722 22473 14738 22507
rect 14772 22473 14784 22507
rect 14722 22439 14784 22473
rect 14722 22405 14738 22439
rect 14772 22405 14784 22439
rect 14722 22371 14784 22405
rect 14722 22337 14738 22371
rect 14772 22337 14784 22371
rect 14722 22303 14784 22337
rect 14722 22269 14738 22303
rect 14772 22269 14784 22303
rect 14722 22235 14784 22269
rect 14722 22201 14738 22235
rect 14772 22201 14784 22235
rect 14722 22167 14784 22201
rect 14722 22133 14738 22167
rect 14772 22133 14784 22167
rect 14722 22099 14784 22133
rect 14722 22065 14738 22099
rect 14772 22065 14784 22099
rect 14722 22031 14784 22065
rect 14722 21997 14738 22031
rect 14772 21997 14784 22031
rect 14722 21963 14784 21997
rect 14722 21929 14738 21963
rect 14772 21929 14784 21963
rect 14722 21895 14784 21929
rect 14722 21861 14738 21895
rect 14772 21861 14784 21895
rect 14722 21827 14784 21861
rect 14722 21793 14738 21827
rect 14772 21793 14784 21827
rect 14722 21759 14784 21793
rect 14722 21725 14738 21759
rect 14772 21725 14784 21759
rect 14722 21691 14784 21725
rect 14722 21657 14738 21691
rect 14772 21657 14784 21691
rect 14722 21623 14784 21657
rect 14722 21589 14738 21623
rect 14772 21589 14784 21623
rect 14722 21555 14784 21589
rect 14722 21521 14738 21555
rect 14772 21521 14784 21555
rect 14722 21487 14784 21521
rect 14722 21453 14738 21487
rect 14772 21453 14784 21487
rect 14722 21419 14784 21453
rect 14722 21385 14738 21419
rect 14772 21385 14784 21419
rect 14722 21351 14784 21385
rect 14722 21317 14738 21351
rect 14772 21317 14784 21351
rect 14722 21283 14784 21317
rect 14722 21249 14738 21283
rect 14772 21249 14784 21283
rect 14722 21215 14784 21249
rect 14722 21181 14738 21215
rect 14772 21181 14784 21215
rect 14722 21150 14784 21181
rect 16650 24009 16712 24040
rect 16650 23975 16662 24009
rect 16696 23975 16712 24009
rect 16650 23941 16712 23975
rect 16650 23907 16662 23941
rect 16696 23907 16712 23941
rect 16650 23873 16712 23907
rect 16650 23839 16662 23873
rect 16696 23839 16712 23873
rect 16650 23805 16712 23839
rect 16650 23771 16662 23805
rect 16696 23771 16712 23805
rect 16650 23737 16712 23771
rect 16650 23703 16662 23737
rect 16696 23703 16712 23737
rect 16650 23669 16712 23703
rect 16650 23635 16662 23669
rect 16696 23635 16712 23669
rect 16650 23601 16712 23635
rect 16650 23567 16662 23601
rect 16696 23567 16712 23601
rect 16650 23533 16712 23567
rect 16650 23499 16662 23533
rect 16696 23499 16712 23533
rect 16650 23465 16712 23499
rect 16650 23431 16662 23465
rect 16696 23431 16712 23465
rect 16650 23397 16712 23431
rect 16650 23363 16662 23397
rect 16696 23363 16712 23397
rect 16650 23329 16712 23363
rect 16650 23295 16662 23329
rect 16696 23295 16712 23329
rect 16650 23261 16712 23295
rect 16650 23227 16662 23261
rect 16696 23227 16712 23261
rect 16650 23193 16712 23227
rect 16650 23159 16662 23193
rect 16696 23159 16712 23193
rect 16650 23125 16712 23159
rect 16650 23091 16662 23125
rect 16696 23091 16712 23125
rect 16650 23057 16712 23091
rect 16650 23023 16662 23057
rect 16696 23023 16712 23057
rect 16650 22989 16712 23023
rect 16650 22955 16662 22989
rect 16696 22955 16712 22989
rect 16650 22921 16712 22955
rect 16650 22887 16662 22921
rect 16696 22887 16712 22921
rect 16650 22853 16712 22887
rect 16650 22819 16662 22853
rect 16696 22819 16712 22853
rect 16650 22785 16712 22819
rect 16650 22751 16662 22785
rect 16696 22751 16712 22785
rect 16650 22717 16712 22751
rect 16650 22683 16662 22717
rect 16696 22683 16712 22717
rect 16650 22649 16712 22683
rect 16650 22615 16662 22649
rect 16696 22615 16712 22649
rect 16650 22581 16712 22615
rect 16650 22547 16662 22581
rect 16696 22547 16712 22581
rect 16650 22513 16712 22547
rect 16650 22479 16662 22513
rect 16696 22479 16712 22513
rect 16650 22445 16712 22479
rect 16650 22411 16662 22445
rect 16696 22411 16712 22445
rect 16650 22377 16712 22411
rect 16650 22343 16662 22377
rect 16696 22343 16712 22377
rect 16650 22309 16712 22343
rect 16650 22275 16662 22309
rect 16696 22275 16712 22309
rect 16650 22241 16712 22275
rect 16650 22207 16662 22241
rect 16696 22207 16712 22241
rect 16650 22173 16712 22207
rect 16650 22139 16662 22173
rect 16696 22139 16712 22173
rect 16650 22105 16712 22139
rect 16650 22071 16662 22105
rect 16696 22071 16712 22105
rect 16650 22040 16712 22071
rect 16742 24009 16808 24040
rect 16742 23975 16758 24009
rect 16792 23975 16808 24009
rect 16742 23941 16808 23975
rect 16742 23907 16758 23941
rect 16792 23907 16808 23941
rect 16742 23873 16808 23907
rect 16742 23839 16758 23873
rect 16792 23839 16808 23873
rect 16742 23805 16808 23839
rect 16742 23771 16758 23805
rect 16792 23771 16808 23805
rect 16742 23737 16808 23771
rect 16742 23703 16758 23737
rect 16792 23703 16808 23737
rect 16742 23669 16808 23703
rect 16742 23635 16758 23669
rect 16792 23635 16808 23669
rect 16742 23601 16808 23635
rect 16742 23567 16758 23601
rect 16792 23567 16808 23601
rect 16742 23533 16808 23567
rect 16742 23499 16758 23533
rect 16792 23499 16808 23533
rect 16742 23465 16808 23499
rect 16742 23431 16758 23465
rect 16792 23431 16808 23465
rect 16742 23397 16808 23431
rect 16742 23363 16758 23397
rect 16792 23363 16808 23397
rect 16742 23329 16808 23363
rect 16742 23295 16758 23329
rect 16792 23295 16808 23329
rect 16742 23261 16808 23295
rect 16742 23227 16758 23261
rect 16792 23227 16808 23261
rect 16742 23193 16808 23227
rect 16742 23159 16758 23193
rect 16792 23159 16808 23193
rect 16742 23125 16808 23159
rect 16742 23091 16758 23125
rect 16792 23091 16808 23125
rect 16742 23057 16808 23091
rect 16742 23023 16758 23057
rect 16792 23023 16808 23057
rect 16742 22989 16808 23023
rect 16742 22955 16758 22989
rect 16792 22955 16808 22989
rect 16742 22921 16808 22955
rect 16742 22887 16758 22921
rect 16792 22887 16808 22921
rect 16742 22853 16808 22887
rect 16742 22819 16758 22853
rect 16792 22819 16808 22853
rect 16742 22785 16808 22819
rect 16742 22751 16758 22785
rect 16792 22751 16808 22785
rect 16742 22717 16808 22751
rect 16742 22683 16758 22717
rect 16792 22683 16808 22717
rect 16742 22649 16808 22683
rect 16742 22615 16758 22649
rect 16792 22615 16808 22649
rect 16742 22581 16808 22615
rect 16742 22547 16758 22581
rect 16792 22547 16808 22581
rect 16742 22513 16808 22547
rect 16742 22479 16758 22513
rect 16792 22479 16808 22513
rect 16742 22445 16808 22479
rect 16742 22411 16758 22445
rect 16792 22411 16808 22445
rect 16742 22377 16808 22411
rect 16742 22343 16758 22377
rect 16792 22343 16808 22377
rect 16742 22309 16808 22343
rect 16742 22275 16758 22309
rect 16792 22275 16808 22309
rect 16742 22241 16808 22275
rect 16742 22207 16758 22241
rect 16792 22207 16808 22241
rect 16742 22173 16808 22207
rect 16742 22139 16758 22173
rect 16792 22139 16808 22173
rect 16742 22105 16808 22139
rect 16742 22071 16758 22105
rect 16792 22071 16808 22105
rect 16742 22040 16808 22071
rect 16838 24009 16904 24040
rect 16838 23975 16854 24009
rect 16888 23975 16904 24009
rect 16838 23941 16904 23975
rect 16838 23907 16854 23941
rect 16888 23907 16904 23941
rect 16838 23873 16904 23907
rect 16838 23839 16854 23873
rect 16888 23839 16904 23873
rect 16838 23805 16904 23839
rect 16838 23771 16854 23805
rect 16888 23771 16904 23805
rect 16838 23737 16904 23771
rect 16838 23703 16854 23737
rect 16888 23703 16904 23737
rect 16838 23669 16904 23703
rect 16838 23635 16854 23669
rect 16888 23635 16904 23669
rect 16838 23601 16904 23635
rect 16838 23567 16854 23601
rect 16888 23567 16904 23601
rect 16838 23533 16904 23567
rect 16838 23499 16854 23533
rect 16888 23499 16904 23533
rect 16838 23465 16904 23499
rect 16838 23431 16854 23465
rect 16888 23431 16904 23465
rect 16838 23397 16904 23431
rect 16838 23363 16854 23397
rect 16888 23363 16904 23397
rect 16838 23329 16904 23363
rect 16838 23295 16854 23329
rect 16888 23295 16904 23329
rect 16838 23261 16904 23295
rect 16838 23227 16854 23261
rect 16888 23227 16904 23261
rect 16838 23193 16904 23227
rect 16838 23159 16854 23193
rect 16888 23159 16904 23193
rect 16838 23125 16904 23159
rect 16838 23091 16854 23125
rect 16888 23091 16904 23125
rect 16838 23057 16904 23091
rect 16838 23023 16854 23057
rect 16888 23023 16904 23057
rect 16838 22989 16904 23023
rect 16838 22955 16854 22989
rect 16888 22955 16904 22989
rect 16838 22921 16904 22955
rect 16838 22887 16854 22921
rect 16888 22887 16904 22921
rect 16838 22853 16904 22887
rect 16838 22819 16854 22853
rect 16888 22819 16904 22853
rect 16838 22785 16904 22819
rect 16838 22751 16854 22785
rect 16888 22751 16904 22785
rect 16838 22717 16904 22751
rect 16838 22683 16854 22717
rect 16888 22683 16904 22717
rect 16838 22649 16904 22683
rect 16838 22615 16854 22649
rect 16888 22615 16904 22649
rect 16838 22581 16904 22615
rect 16838 22547 16854 22581
rect 16888 22547 16904 22581
rect 16838 22513 16904 22547
rect 16838 22479 16854 22513
rect 16888 22479 16904 22513
rect 16838 22445 16904 22479
rect 16838 22411 16854 22445
rect 16888 22411 16904 22445
rect 16838 22377 16904 22411
rect 16838 22343 16854 22377
rect 16888 22343 16904 22377
rect 16838 22309 16904 22343
rect 16838 22275 16854 22309
rect 16888 22275 16904 22309
rect 16838 22241 16904 22275
rect 16838 22207 16854 22241
rect 16888 22207 16904 22241
rect 16838 22173 16904 22207
rect 16838 22139 16854 22173
rect 16888 22139 16904 22173
rect 16838 22105 16904 22139
rect 16838 22071 16854 22105
rect 16888 22071 16904 22105
rect 16838 22040 16904 22071
rect 16934 24009 17000 24040
rect 16934 23975 16950 24009
rect 16984 23975 17000 24009
rect 16934 23941 17000 23975
rect 16934 23907 16950 23941
rect 16984 23907 17000 23941
rect 16934 23873 17000 23907
rect 16934 23839 16950 23873
rect 16984 23839 17000 23873
rect 16934 23805 17000 23839
rect 16934 23771 16950 23805
rect 16984 23771 17000 23805
rect 16934 23737 17000 23771
rect 16934 23703 16950 23737
rect 16984 23703 17000 23737
rect 16934 23669 17000 23703
rect 16934 23635 16950 23669
rect 16984 23635 17000 23669
rect 16934 23601 17000 23635
rect 16934 23567 16950 23601
rect 16984 23567 17000 23601
rect 16934 23533 17000 23567
rect 16934 23499 16950 23533
rect 16984 23499 17000 23533
rect 16934 23465 17000 23499
rect 16934 23431 16950 23465
rect 16984 23431 17000 23465
rect 16934 23397 17000 23431
rect 16934 23363 16950 23397
rect 16984 23363 17000 23397
rect 16934 23329 17000 23363
rect 16934 23295 16950 23329
rect 16984 23295 17000 23329
rect 16934 23261 17000 23295
rect 16934 23227 16950 23261
rect 16984 23227 17000 23261
rect 16934 23193 17000 23227
rect 16934 23159 16950 23193
rect 16984 23159 17000 23193
rect 16934 23125 17000 23159
rect 16934 23091 16950 23125
rect 16984 23091 17000 23125
rect 16934 23057 17000 23091
rect 16934 23023 16950 23057
rect 16984 23023 17000 23057
rect 16934 22989 17000 23023
rect 16934 22955 16950 22989
rect 16984 22955 17000 22989
rect 16934 22921 17000 22955
rect 16934 22887 16950 22921
rect 16984 22887 17000 22921
rect 16934 22853 17000 22887
rect 16934 22819 16950 22853
rect 16984 22819 17000 22853
rect 16934 22785 17000 22819
rect 16934 22751 16950 22785
rect 16984 22751 17000 22785
rect 16934 22717 17000 22751
rect 16934 22683 16950 22717
rect 16984 22683 17000 22717
rect 16934 22649 17000 22683
rect 16934 22615 16950 22649
rect 16984 22615 17000 22649
rect 16934 22581 17000 22615
rect 16934 22547 16950 22581
rect 16984 22547 17000 22581
rect 16934 22513 17000 22547
rect 16934 22479 16950 22513
rect 16984 22479 17000 22513
rect 16934 22445 17000 22479
rect 16934 22411 16950 22445
rect 16984 22411 17000 22445
rect 16934 22377 17000 22411
rect 16934 22343 16950 22377
rect 16984 22343 17000 22377
rect 16934 22309 17000 22343
rect 16934 22275 16950 22309
rect 16984 22275 17000 22309
rect 16934 22241 17000 22275
rect 16934 22207 16950 22241
rect 16984 22207 17000 22241
rect 16934 22173 17000 22207
rect 16934 22139 16950 22173
rect 16984 22139 17000 22173
rect 16934 22105 17000 22139
rect 16934 22071 16950 22105
rect 16984 22071 17000 22105
rect 16934 22040 17000 22071
rect 17030 24009 17096 24040
rect 17030 23975 17046 24009
rect 17080 23975 17096 24009
rect 17030 23941 17096 23975
rect 17030 23907 17046 23941
rect 17080 23907 17096 23941
rect 17030 23873 17096 23907
rect 17030 23839 17046 23873
rect 17080 23839 17096 23873
rect 17030 23805 17096 23839
rect 17030 23771 17046 23805
rect 17080 23771 17096 23805
rect 17030 23737 17096 23771
rect 17030 23703 17046 23737
rect 17080 23703 17096 23737
rect 17030 23669 17096 23703
rect 17030 23635 17046 23669
rect 17080 23635 17096 23669
rect 17030 23601 17096 23635
rect 17030 23567 17046 23601
rect 17080 23567 17096 23601
rect 17030 23533 17096 23567
rect 17030 23499 17046 23533
rect 17080 23499 17096 23533
rect 17030 23465 17096 23499
rect 17030 23431 17046 23465
rect 17080 23431 17096 23465
rect 17030 23397 17096 23431
rect 17030 23363 17046 23397
rect 17080 23363 17096 23397
rect 17030 23329 17096 23363
rect 17030 23295 17046 23329
rect 17080 23295 17096 23329
rect 17030 23261 17096 23295
rect 17030 23227 17046 23261
rect 17080 23227 17096 23261
rect 17030 23193 17096 23227
rect 17030 23159 17046 23193
rect 17080 23159 17096 23193
rect 17030 23125 17096 23159
rect 17030 23091 17046 23125
rect 17080 23091 17096 23125
rect 17030 23057 17096 23091
rect 17030 23023 17046 23057
rect 17080 23023 17096 23057
rect 17030 22989 17096 23023
rect 17030 22955 17046 22989
rect 17080 22955 17096 22989
rect 17030 22921 17096 22955
rect 17030 22887 17046 22921
rect 17080 22887 17096 22921
rect 17030 22853 17096 22887
rect 17030 22819 17046 22853
rect 17080 22819 17096 22853
rect 17030 22785 17096 22819
rect 17030 22751 17046 22785
rect 17080 22751 17096 22785
rect 17030 22717 17096 22751
rect 17030 22683 17046 22717
rect 17080 22683 17096 22717
rect 17030 22649 17096 22683
rect 17030 22615 17046 22649
rect 17080 22615 17096 22649
rect 17030 22581 17096 22615
rect 17030 22547 17046 22581
rect 17080 22547 17096 22581
rect 17030 22513 17096 22547
rect 17030 22479 17046 22513
rect 17080 22479 17096 22513
rect 17030 22445 17096 22479
rect 17030 22411 17046 22445
rect 17080 22411 17096 22445
rect 17030 22377 17096 22411
rect 17030 22343 17046 22377
rect 17080 22343 17096 22377
rect 17030 22309 17096 22343
rect 17030 22275 17046 22309
rect 17080 22275 17096 22309
rect 17030 22241 17096 22275
rect 17030 22207 17046 22241
rect 17080 22207 17096 22241
rect 17030 22173 17096 22207
rect 17030 22139 17046 22173
rect 17080 22139 17096 22173
rect 17030 22105 17096 22139
rect 17030 22071 17046 22105
rect 17080 22071 17096 22105
rect 17030 22040 17096 22071
rect 17126 24009 17192 24040
rect 17126 23975 17142 24009
rect 17176 23975 17192 24009
rect 17126 23941 17192 23975
rect 17126 23907 17142 23941
rect 17176 23907 17192 23941
rect 17126 23873 17192 23907
rect 17126 23839 17142 23873
rect 17176 23839 17192 23873
rect 17126 23805 17192 23839
rect 17126 23771 17142 23805
rect 17176 23771 17192 23805
rect 17126 23737 17192 23771
rect 17126 23703 17142 23737
rect 17176 23703 17192 23737
rect 17126 23669 17192 23703
rect 17126 23635 17142 23669
rect 17176 23635 17192 23669
rect 17126 23601 17192 23635
rect 17126 23567 17142 23601
rect 17176 23567 17192 23601
rect 17126 23533 17192 23567
rect 17126 23499 17142 23533
rect 17176 23499 17192 23533
rect 17126 23465 17192 23499
rect 17126 23431 17142 23465
rect 17176 23431 17192 23465
rect 17126 23397 17192 23431
rect 17126 23363 17142 23397
rect 17176 23363 17192 23397
rect 17126 23329 17192 23363
rect 17126 23295 17142 23329
rect 17176 23295 17192 23329
rect 17126 23261 17192 23295
rect 17126 23227 17142 23261
rect 17176 23227 17192 23261
rect 17126 23193 17192 23227
rect 17126 23159 17142 23193
rect 17176 23159 17192 23193
rect 17126 23125 17192 23159
rect 17126 23091 17142 23125
rect 17176 23091 17192 23125
rect 17126 23057 17192 23091
rect 17126 23023 17142 23057
rect 17176 23023 17192 23057
rect 17126 22989 17192 23023
rect 17126 22955 17142 22989
rect 17176 22955 17192 22989
rect 17126 22921 17192 22955
rect 17126 22887 17142 22921
rect 17176 22887 17192 22921
rect 17126 22853 17192 22887
rect 17126 22819 17142 22853
rect 17176 22819 17192 22853
rect 17126 22785 17192 22819
rect 17126 22751 17142 22785
rect 17176 22751 17192 22785
rect 17126 22717 17192 22751
rect 17126 22683 17142 22717
rect 17176 22683 17192 22717
rect 17126 22649 17192 22683
rect 17126 22615 17142 22649
rect 17176 22615 17192 22649
rect 17126 22581 17192 22615
rect 17126 22547 17142 22581
rect 17176 22547 17192 22581
rect 17126 22513 17192 22547
rect 17126 22479 17142 22513
rect 17176 22479 17192 22513
rect 17126 22445 17192 22479
rect 17126 22411 17142 22445
rect 17176 22411 17192 22445
rect 17126 22377 17192 22411
rect 17126 22343 17142 22377
rect 17176 22343 17192 22377
rect 17126 22309 17192 22343
rect 17126 22275 17142 22309
rect 17176 22275 17192 22309
rect 17126 22241 17192 22275
rect 17126 22207 17142 22241
rect 17176 22207 17192 22241
rect 17126 22173 17192 22207
rect 17126 22139 17142 22173
rect 17176 22139 17192 22173
rect 17126 22105 17192 22139
rect 17126 22071 17142 22105
rect 17176 22071 17192 22105
rect 17126 22040 17192 22071
rect 17222 24009 17288 24040
rect 17222 23975 17238 24009
rect 17272 23975 17288 24009
rect 17222 23941 17288 23975
rect 17222 23907 17238 23941
rect 17272 23907 17288 23941
rect 17222 23873 17288 23907
rect 17222 23839 17238 23873
rect 17272 23839 17288 23873
rect 17222 23805 17288 23839
rect 17222 23771 17238 23805
rect 17272 23771 17288 23805
rect 17222 23737 17288 23771
rect 17222 23703 17238 23737
rect 17272 23703 17288 23737
rect 17222 23669 17288 23703
rect 17222 23635 17238 23669
rect 17272 23635 17288 23669
rect 17222 23601 17288 23635
rect 17222 23567 17238 23601
rect 17272 23567 17288 23601
rect 17222 23533 17288 23567
rect 17222 23499 17238 23533
rect 17272 23499 17288 23533
rect 17222 23465 17288 23499
rect 17222 23431 17238 23465
rect 17272 23431 17288 23465
rect 17222 23397 17288 23431
rect 17222 23363 17238 23397
rect 17272 23363 17288 23397
rect 17222 23329 17288 23363
rect 17222 23295 17238 23329
rect 17272 23295 17288 23329
rect 17222 23261 17288 23295
rect 17222 23227 17238 23261
rect 17272 23227 17288 23261
rect 17222 23193 17288 23227
rect 17222 23159 17238 23193
rect 17272 23159 17288 23193
rect 17222 23125 17288 23159
rect 17222 23091 17238 23125
rect 17272 23091 17288 23125
rect 17222 23057 17288 23091
rect 17222 23023 17238 23057
rect 17272 23023 17288 23057
rect 17222 22989 17288 23023
rect 17222 22955 17238 22989
rect 17272 22955 17288 22989
rect 17222 22921 17288 22955
rect 17222 22887 17238 22921
rect 17272 22887 17288 22921
rect 17222 22853 17288 22887
rect 17222 22819 17238 22853
rect 17272 22819 17288 22853
rect 17222 22785 17288 22819
rect 17222 22751 17238 22785
rect 17272 22751 17288 22785
rect 17222 22717 17288 22751
rect 17222 22683 17238 22717
rect 17272 22683 17288 22717
rect 17222 22649 17288 22683
rect 17222 22615 17238 22649
rect 17272 22615 17288 22649
rect 17222 22581 17288 22615
rect 17222 22547 17238 22581
rect 17272 22547 17288 22581
rect 17222 22513 17288 22547
rect 17222 22479 17238 22513
rect 17272 22479 17288 22513
rect 17222 22445 17288 22479
rect 17222 22411 17238 22445
rect 17272 22411 17288 22445
rect 17222 22377 17288 22411
rect 17222 22343 17238 22377
rect 17272 22343 17288 22377
rect 17222 22309 17288 22343
rect 17222 22275 17238 22309
rect 17272 22275 17288 22309
rect 17222 22241 17288 22275
rect 17222 22207 17238 22241
rect 17272 22207 17288 22241
rect 17222 22173 17288 22207
rect 17222 22139 17238 22173
rect 17272 22139 17288 22173
rect 17222 22105 17288 22139
rect 17222 22071 17238 22105
rect 17272 22071 17288 22105
rect 17222 22040 17288 22071
rect 17318 24009 17384 24040
rect 17318 23975 17334 24009
rect 17368 23975 17384 24009
rect 17318 23941 17384 23975
rect 17318 23907 17334 23941
rect 17368 23907 17384 23941
rect 17318 23873 17384 23907
rect 17318 23839 17334 23873
rect 17368 23839 17384 23873
rect 17318 23805 17384 23839
rect 17318 23771 17334 23805
rect 17368 23771 17384 23805
rect 17318 23737 17384 23771
rect 17318 23703 17334 23737
rect 17368 23703 17384 23737
rect 17318 23669 17384 23703
rect 17318 23635 17334 23669
rect 17368 23635 17384 23669
rect 17318 23601 17384 23635
rect 17318 23567 17334 23601
rect 17368 23567 17384 23601
rect 17318 23533 17384 23567
rect 17318 23499 17334 23533
rect 17368 23499 17384 23533
rect 17318 23465 17384 23499
rect 17318 23431 17334 23465
rect 17368 23431 17384 23465
rect 17318 23397 17384 23431
rect 17318 23363 17334 23397
rect 17368 23363 17384 23397
rect 17318 23329 17384 23363
rect 17318 23295 17334 23329
rect 17368 23295 17384 23329
rect 17318 23261 17384 23295
rect 17318 23227 17334 23261
rect 17368 23227 17384 23261
rect 17318 23193 17384 23227
rect 17318 23159 17334 23193
rect 17368 23159 17384 23193
rect 17318 23125 17384 23159
rect 17318 23091 17334 23125
rect 17368 23091 17384 23125
rect 17318 23057 17384 23091
rect 17318 23023 17334 23057
rect 17368 23023 17384 23057
rect 17318 22989 17384 23023
rect 17318 22955 17334 22989
rect 17368 22955 17384 22989
rect 17318 22921 17384 22955
rect 17318 22887 17334 22921
rect 17368 22887 17384 22921
rect 17318 22853 17384 22887
rect 17318 22819 17334 22853
rect 17368 22819 17384 22853
rect 17318 22785 17384 22819
rect 17318 22751 17334 22785
rect 17368 22751 17384 22785
rect 17318 22717 17384 22751
rect 17318 22683 17334 22717
rect 17368 22683 17384 22717
rect 17318 22649 17384 22683
rect 17318 22615 17334 22649
rect 17368 22615 17384 22649
rect 17318 22581 17384 22615
rect 17318 22547 17334 22581
rect 17368 22547 17384 22581
rect 17318 22513 17384 22547
rect 17318 22479 17334 22513
rect 17368 22479 17384 22513
rect 17318 22445 17384 22479
rect 17318 22411 17334 22445
rect 17368 22411 17384 22445
rect 17318 22377 17384 22411
rect 17318 22343 17334 22377
rect 17368 22343 17384 22377
rect 17318 22309 17384 22343
rect 17318 22275 17334 22309
rect 17368 22275 17384 22309
rect 17318 22241 17384 22275
rect 17318 22207 17334 22241
rect 17368 22207 17384 22241
rect 17318 22173 17384 22207
rect 17318 22139 17334 22173
rect 17368 22139 17384 22173
rect 17318 22105 17384 22139
rect 17318 22071 17334 22105
rect 17368 22071 17384 22105
rect 17318 22040 17384 22071
rect 17414 24009 17480 24040
rect 17414 23975 17430 24009
rect 17464 23975 17480 24009
rect 17414 23941 17480 23975
rect 17414 23907 17430 23941
rect 17464 23907 17480 23941
rect 17414 23873 17480 23907
rect 17414 23839 17430 23873
rect 17464 23839 17480 23873
rect 17414 23805 17480 23839
rect 17414 23771 17430 23805
rect 17464 23771 17480 23805
rect 17414 23737 17480 23771
rect 17414 23703 17430 23737
rect 17464 23703 17480 23737
rect 17414 23669 17480 23703
rect 17414 23635 17430 23669
rect 17464 23635 17480 23669
rect 17414 23601 17480 23635
rect 17414 23567 17430 23601
rect 17464 23567 17480 23601
rect 17414 23533 17480 23567
rect 17414 23499 17430 23533
rect 17464 23499 17480 23533
rect 17414 23465 17480 23499
rect 17414 23431 17430 23465
rect 17464 23431 17480 23465
rect 17414 23397 17480 23431
rect 17414 23363 17430 23397
rect 17464 23363 17480 23397
rect 17414 23329 17480 23363
rect 17414 23295 17430 23329
rect 17464 23295 17480 23329
rect 17414 23261 17480 23295
rect 17414 23227 17430 23261
rect 17464 23227 17480 23261
rect 17414 23193 17480 23227
rect 17414 23159 17430 23193
rect 17464 23159 17480 23193
rect 17414 23125 17480 23159
rect 17414 23091 17430 23125
rect 17464 23091 17480 23125
rect 17414 23057 17480 23091
rect 17414 23023 17430 23057
rect 17464 23023 17480 23057
rect 17414 22989 17480 23023
rect 17414 22955 17430 22989
rect 17464 22955 17480 22989
rect 17414 22921 17480 22955
rect 17414 22887 17430 22921
rect 17464 22887 17480 22921
rect 17414 22853 17480 22887
rect 17414 22819 17430 22853
rect 17464 22819 17480 22853
rect 17414 22785 17480 22819
rect 17414 22751 17430 22785
rect 17464 22751 17480 22785
rect 17414 22717 17480 22751
rect 17414 22683 17430 22717
rect 17464 22683 17480 22717
rect 17414 22649 17480 22683
rect 17414 22615 17430 22649
rect 17464 22615 17480 22649
rect 17414 22581 17480 22615
rect 17414 22547 17430 22581
rect 17464 22547 17480 22581
rect 17414 22513 17480 22547
rect 17414 22479 17430 22513
rect 17464 22479 17480 22513
rect 17414 22445 17480 22479
rect 17414 22411 17430 22445
rect 17464 22411 17480 22445
rect 17414 22377 17480 22411
rect 17414 22343 17430 22377
rect 17464 22343 17480 22377
rect 17414 22309 17480 22343
rect 17414 22275 17430 22309
rect 17464 22275 17480 22309
rect 17414 22241 17480 22275
rect 17414 22207 17430 22241
rect 17464 22207 17480 22241
rect 17414 22173 17480 22207
rect 17414 22139 17430 22173
rect 17464 22139 17480 22173
rect 17414 22105 17480 22139
rect 17414 22071 17430 22105
rect 17464 22071 17480 22105
rect 17414 22040 17480 22071
rect 17510 24009 17576 24040
rect 17510 23975 17526 24009
rect 17560 23975 17576 24009
rect 17510 23941 17576 23975
rect 17510 23907 17526 23941
rect 17560 23907 17576 23941
rect 17510 23873 17576 23907
rect 17510 23839 17526 23873
rect 17560 23839 17576 23873
rect 17510 23805 17576 23839
rect 17510 23771 17526 23805
rect 17560 23771 17576 23805
rect 17510 23737 17576 23771
rect 17510 23703 17526 23737
rect 17560 23703 17576 23737
rect 17510 23669 17576 23703
rect 17510 23635 17526 23669
rect 17560 23635 17576 23669
rect 17510 23601 17576 23635
rect 17510 23567 17526 23601
rect 17560 23567 17576 23601
rect 17510 23533 17576 23567
rect 17510 23499 17526 23533
rect 17560 23499 17576 23533
rect 17510 23465 17576 23499
rect 17510 23431 17526 23465
rect 17560 23431 17576 23465
rect 17510 23397 17576 23431
rect 17510 23363 17526 23397
rect 17560 23363 17576 23397
rect 17510 23329 17576 23363
rect 17510 23295 17526 23329
rect 17560 23295 17576 23329
rect 17510 23261 17576 23295
rect 17510 23227 17526 23261
rect 17560 23227 17576 23261
rect 17510 23193 17576 23227
rect 17510 23159 17526 23193
rect 17560 23159 17576 23193
rect 17510 23125 17576 23159
rect 17510 23091 17526 23125
rect 17560 23091 17576 23125
rect 17510 23057 17576 23091
rect 17510 23023 17526 23057
rect 17560 23023 17576 23057
rect 17510 22989 17576 23023
rect 17510 22955 17526 22989
rect 17560 22955 17576 22989
rect 17510 22921 17576 22955
rect 17510 22887 17526 22921
rect 17560 22887 17576 22921
rect 17510 22853 17576 22887
rect 17510 22819 17526 22853
rect 17560 22819 17576 22853
rect 17510 22785 17576 22819
rect 17510 22751 17526 22785
rect 17560 22751 17576 22785
rect 17510 22717 17576 22751
rect 17510 22683 17526 22717
rect 17560 22683 17576 22717
rect 17510 22649 17576 22683
rect 17510 22615 17526 22649
rect 17560 22615 17576 22649
rect 17510 22581 17576 22615
rect 17510 22547 17526 22581
rect 17560 22547 17576 22581
rect 17510 22513 17576 22547
rect 17510 22479 17526 22513
rect 17560 22479 17576 22513
rect 17510 22445 17576 22479
rect 17510 22411 17526 22445
rect 17560 22411 17576 22445
rect 17510 22377 17576 22411
rect 17510 22343 17526 22377
rect 17560 22343 17576 22377
rect 17510 22309 17576 22343
rect 17510 22275 17526 22309
rect 17560 22275 17576 22309
rect 17510 22241 17576 22275
rect 17510 22207 17526 22241
rect 17560 22207 17576 22241
rect 17510 22173 17576 22207
rect 17510 22139 17526 22173
rect 17560 22139 17576 22173
rect 17510 22105 17576 22139
rect 17510 22071 17526 22105
rect 17560 22071 17576 22105
rect 17510 22040 17576 22071
rect 17606 24009 17668 24040
rect 17606 23975 17622 24009
rect 17656 23975 17668 24009
rect 17606 23941 17668 23975
rect 17606 23907 17622 23941
rect 17656 23907 17668 23941
rect 17606 23873 17668 23907
rect 17606 23839 17622 23873
rect 17656 23839 17668 23873
rect 17606 23805 17668 23839
rect 17606 23771 17622 23805
rect 17656 23771 17668 23805
rect 17606 23737 17668 23771
rect 17606 23703 17622 23737
rect 17656 23703 17668 23737
rect 17606 23669 17668 23703
rect 17606 23635 17622 23669
rect 17656 23635 17668 23669
rect 17606 23601 17668 23635
rect 17606 23567 17622 23601
rect 17656 23567 17668 23601
rect 17606 23533 17668 23567
rect 17606 23499 17622 23533
rect 17656 23499 17668 23533
rect 17606 23465 17668 23499
rect 17606 23431 17622 23465
rect 17656 23431 17668 23465
rect 17606 23397 17668 23431
rect 17606 23363 17622 23397
rect 17656 23363 17668 23397
rect 17606 23329 17668 23363
rect 17606 23295 17622 23329
rect 17656 23295 17668 23329
rect 17606 23261 17668 23295
rect 17606 23227 17622 23261
rect 17656 23227 17668 23261
rect 17606 23193 17668 23227
rect 17606 23159 17622 23193
rect 17656 23159 17668 23193
rect 17606 23125 17668 23159
rect 17606 23091 17622 23125
rect 17656 23091 17668 23125
rect 17606 23057 17668 23091
rect 17606 23023 17622 23057
rect 17656 23023 17668 23057
rect 17606 22989 17668 23023
rect 17606 22955 17622 22989
rect 17656 22955 17668 22989
rect 17606 22921 17668 22955
rect 17606 22887 17622 22921
rect 17656 22887 17668 22921
rect 17606 22853 17668 22887
rect 17606 22819 17622 22853
rect 17656 22819 17668 22853
rect 17606 22785 17668 22819
rect 17606 22751 17622 22785
rect 17656 22751 17668 22785
rect 17606 22717 17668 22751
rect 17606 22683 17622 22717
rect 17656 22683 17668 22717
rect 17606 22649 17668 22683
rect 17606 22615 17622 22649
rect 17656 22615 17668 22649
rect 17606 22581 17668 22615
rect 17606 22547 17622 22581
rect 17656 22547 17668 22581
rect 17606 22513 17668 22547
rect 17606 22479 17622 22513
rect 17656 22479 17668 22513
rect 17606 22445 17668 22479
rect 17606 22411 17622 22445
rect 17656 22411 17668 22445
rect 17606 22377 17668 22411
rect 17606 22343 17622 22377
rect 17656 22343 17668 22377
rect 17606 22309 17668 22343
rect 17606 22275 17622 22309
rect 17656 22275 17668 22309
rect 17606 22241 17668 22275
rect 17606 22207 17622 22241
rect 17656 22207 17668 22241
rect 17606 22173 17668 22207
rect 17606 22139 17622 22173
rect 17656 22139 17668 22173
rect 17606 22105 17668 22139
rect 17606 22071 17622 22105
rect 17656 22071 17668 22105
rect 17606 22040 17668 22071
rect 14818 20432 14880 20446
rect 14818 20398 14830 20432
rect 14864 20398 14880 20432
rect 14818 20364 14880 20398
rect 14818 20330 14830 20364
rect 14864 20330 14880 20364
rect 14818 20296 14880 20330
rect 14818 20262 14830 20296
rect 14864 20262 14880 20296
rect 14818 20228 14880 20262
rect 14818 20194 14830 20228
rect 14864 20194 14880 20228
rect 14818 20160 14880 20194
rect 14818 20126 14830 20160
rect 14864 20126 14880 20160
rect 14818 20092 14880 20126
rect 14818 20058 14830 20092
rect 14864 20058 14880 20092
rect 14818 20024 14880 20058
rect 14818 19990 14830 20024
rect 14864 19990 14880 20024
rect 14818 19956 14880 19990
rect 14818 19922 14830 19956
rect 14864 19922 14880 19956
rect 14818 19888 14880 19922
rect 14818 19854 14830 19888
rect 14864 19854 14880 19888
rect 14818 19820 14880 19854
rect 14818 19786 14830 19820
rect 14864 19786 14880 19820
rect 14818 19752 14880 19786
rect 14818 19718 14830 19752
rect 14864 19718 14880 19752
rect 14818 19684 14880 19718
rect 14818 19650 14830 19684
rect 14864 19650 14880 19684
rect 14818 19616 14880 19650
rect 14818 19582 14830 19616
rect 14864 19582 14880 19616
rect 14818 19548 14880 19582
rect 14818 19514 14830 19548
rect 14864 19514 14880 19548
rect 14818 19480 14880 19514
rect 14818 19446 14830 19480
rect 14864 19446 14880 19480
rect 14818 19412 14880 19446
rect 14818 19378 14830 19412
rect 14864 19378 14880 19412
rect 14818 19344 14880 19378
rect 14818 19310 14830 19344
rect 14864 19310 14880 19344
rect 14818 19276 14880 19310
rect 14818 19242 14830 19276
rect 14864 19242 14880 19276
rect 14818 19208 14880 19242
rect 14818 19174 14830 19208
rect 14864 19174 14880 19208
rect 14818 19160 14880 19174
rect 14910 20432 14976 20446
rect 14910 20398 14926 20432
rect 14960 20398 14976 20432
rect 14910 20364 14976 20398
rect 14910 20330 14926 20364
rect 14960 20330 14976 20364
rect 14910 20296 14976 20330
rect 14910 20262 14926 20296
rect 14960 20262 14976 20296
rect 14910 20228 14976 20262
rect 14910 20194 14926 20228
rect 14960 20194 14976 20228
rect 14910 20160 14976 20194
rect 14910 20126 14926 20160
rect 14960 20126 14976 20160
rect 14910 20092 14976 20126
rect 14910 20058 14926 20092
rect 14960 20058 14976 20092
rect 14910 20024 14976 20058
rect 14910 19990 14926 20024
rect 14960 19990 14976 20024
rect 14910 19956 14976 19990
rect 14910 19922 14926 19956
rect 14960 19922 14976 19956
rect 14910 19888 14976 19922
rect 14910 19854 14926 19888
rect 14960 19854 14976 19888
rect 14910 19820 14976 19854
rect 14910 19786 14926 19820
rect 14960 19786 14976 19820
rect 14910 19752 14976 19786
rect 14910 19718 14926 19752
rect 14960 19718 14976 19752
rect 14910 19684 14976 19718
rect 14910 19650 14926 19684
rect 14960 19650 14976 19684
rect 14910 19616 14976 19650
rect 14910 19582 14926 19616
rect 14960 19582 14976 19616
rect 14910 19548 14976 19582
rect 14910 19514 14926 19548
rect 14960 19514 14976 19548
rect 14910 19480 14976 19514
rect 14910 19446 14926 19480
rect 14960 19446 14976 19480
rect 14910 19412 14976 19446
rect 14910 19378 14926 19412
rect 14960 19378 14976 19412
rect 14910 19344 14976 19378
rect 14910 19310 14926 19344
rect 14960 19310 14976 19344
rect 14910 19276 14976 19310
rect 14910 19242 14926 19276
rect 14960 19242 14976 19276
rect 14910 19208 14976 19242
rect 14910 19174 14926 19208
rect 14960 19174 14976 19208
rect 14910 19160 14976 19174
rect 15006 20432 15072 20446
rect 15006 20398 15022 20432
rect 15056 20398 15072 20432
rect 15006 20364 15072 20398
rect 15006 20330 15022 20364
rect 15056 20330 15072 20364
rect 15006 20296 15072 20330
rect 15006 20262 15022 20296
rect 15056 20262 15072 20296
rect 15006 20228 15072 20262
rect 15006 20194 15022 20228
rect 15056 20194 15072 20228
rect 15006 20160 15072 20194
rect 15006 20126 15022 20160
rect 15056 20126 15072 20160
rect 15006 20092 15072 20126
rect 15006 20058 15022 20092
rect 15056 20058 15072 20092
rect 15006 20024 15072 20058
rect 15006 19990 15022 20024
rect 15056 19990 15072 20024
rect 15006 19956 15072 19990
rect 15006 19922 15022 19956
rect 15056 19922 15072 19956
rect 15006 19888 15072 19922
rect 15006 19854 15022 19888
rect 15056 19854 15072 19888
rect 15006 19820 15072 19854
rect 15006 19786 15022 19820
rect 15056 19786 15072 19820
rect 15006 19752 15072 19786
rect 15006 19718 15022 19752
rect 15056 19718 15072 19752
rect 15006 19684 15072 19718
rect 15006 19650 15022 19684
rect 15056 19650 15072 19684
rect 15006 19616 15072 19650
rect 15006 19582 15022 19616
rect 15056 19582 15072 19616
rect 15006 19548 15072 19582
rect 15006 19514 15022 19548
rect 15056 19514 15072 19548
rect 15006 19480 15072 19514
rect 15006 19446 15022 19480
rect 15056 19446 15072 19480
rect 15006 19412 15072 19446
rect 15006 19378 15022 19412
rect 15056 19378 15072 19412
rect 15006 19344 15072 19378
rect 15006 19310 15022 19344
rect 15056 19310 15072 19344
rect 15006 19276 15072 19310
rect 15006 19242 15022 19276
rect 15056 19242 15072 19276
rect 15006 19208 15072 19242
rect 15006 19174 15022 19208
rect 15056 19174 15072 19208
rect 15006 19160 15072 19174
rect 15102 20432 15168 20446
rect 15102 20398 15118 20432
rect 15152 20398 15168 20432
rect 15102 20364 15168 20398
rect 15102 20330 15118 20364
rect 15152 20330 15168 20364
rect 15102 20296 15168 20330
rect 15102 20262 15118 20296
rect 15152 20262 15168 20296
rect 15102 20228 15168 20262
rect 15102 20194 15118 20228
rect 15152 20194 15168 20228
rect 15102 20160 15168 20194
rect 15102 20126 15118 20160
rect 15152 20126 15168 20160
rect 15102 20092 15168 20126
rect 15102 20058 15118 20092
rect 15152 20058 15168 20092
rect 15102 20024 15168 20058
rect 15102 19990 15118 20024
rect 15152 19990 15168 20024
rect 15102 19956 15168 19990
rect 15102 19922 15118 19956
rect 15152 19922 15168 19956
rect 15102 19888 15168 19922
rect 15102 19854 15118 19888
rect 15152 19854 15168 19888
rect 15102 19820 15168 19854
rect 15102 19786 15118 19820
rect 15152 19786 15168 19820
rect 15102 19752 15168 19786
rect 15102 19718 15118 19752
rect 15152 19718 15168 19752
rect 15102 19684 15168 19718
rect 15102 19650 15118 19684
rect 15152 19650 15168 19684
rect 15102 19616 15168 19650
rect 15102 19582 15118 19616
rect 15152 19582 15168 19616
rect 15102 19548 15168 19582
rect 15102 19514 15118 19548
rect 15152 19514 15168 19548
rect 15102 19480 15168 19514
rect 15102 19446 15118 19480
rect 15152 19446 15168 19480
rect 15102 19412 15168 19446
rect 15102 19378 15118 19412
rect 15152 19378 15168 19412
rect 15102 19344 15168 19378
rect 15102 19310 15118 19344
rect 15152 19310 15168 19344
rect 15102 19276 15168 19310
rect 15102 19242 15118 19276
rect 15152 19242 15168 19276
rect 15102 19208 15168 19242
rect 15102 19174 15118 19208
rect 15152 19174 15168 19208
rect 15102 19160 15168 19174
rect 15198 20432 15264 20446
rect 15198 20398 15214 20432
rect 15248 20398 15264 20432
rect 15198 20364 15264 20398
rect 15198 20330 15214 20364
rect 15248 20330 15264 20364
rect 15198 20296 15264 20330
rect 15198 20262 15214 20296
rect 15248 20262 15264 20296
rect 15198 20228 15264 20262
rect 15198 20194 15214 20228
rect 15248 20194 15264 20228
rect 15198 20160 15264 20194
rect 15198 20126 15214 20160
rect 15248 20126 15264 20160
rect 15198 20092 15264 20126
rect 15198 20058 15214 20092
rect 15248 20058 15264 20092
rect 15198 20024 15264 20058
rect 15198 19990 15214 20024
rect 15248 19990 15264 20024
rect 15198 19956 15264 19990
rect 15198 19922 15214 19956
rect 15248 19922 15264 19956
rect 15198 19888 15264 19922
rect 15198 19854 15214 19888
rect 15248 19854 15264 19888
rect 15198 19820 15264 19854
rect 15198 19786 15214 19820
rect 15248 19786 15264 19820
rect 15198 19752 15264 19786
rect 15198 19718 15214 19752
rect 15248 19718 15264 19752
rect 15198 19684 15264 19718
rect 15198 19650 15214 19684
rect 15248 19650 15264 19684
rect 15198 19616 15264 19650
rect 15198 19582 15214 19616
rect 15248 19582 15264 19616
rect 15198 19548 15264 19582
rect 15198 19514 15214 19548
rect 15248 19514 15264 19548
rect 15198 19480 15264 19514
rect 15198 19446 15214 19480
rect 15248 19446 15264 19480
rect 15198 19412 15264 19446
rect 15198 19378 15214 19412
rect 15248 19378 15264 19412
rect 15198 19344 15264 19378
rect 15198 19310 15214 19344
rect 15248 19310 15264 19344
rect 15198 19276 15264 19310
rect 15198 19242 15214 19276
rect 15248 19242 15264 19276
rect 15198 19208 15264 19242
rect 15198 19174 15214 19208
rect 15248 19174 15264 19208
rect 15198 19160 15264 19174
rect 15294 20432 15360 20446
rect 15294 20398 15310 20432
rect 15344 20398 15360 20432
rect 15294 20364 15360 20398
rect 15294 20330 15310 20364
rect 15344 20330 15360 20364
rect 15294 20296 15360 20330
rect 15294 20262 15310 20296
rect 15344 20262 15360 20296
rect 15294 20228 15360 20262
rect 15294 20194 15310 20228
rect 15344 20194 15360 20228
rect 15294 20160 15360 20194
rect 15294 20126 15310 20160
rect 15344 20126 15360 20160
rect 15294 20092 15360 20126
rect 15294 20058 15310 20092
rect 15344 20058 15360 20092
rect 15294 20024 15360 20058
rect 15294 19990 15310 20024
rect 15344 19990 15360 20024
rect 15294 19956 15360 19990
rect 15294 19922 15310 19956
rect 15344 19922 15360 19956
rect 15294 19888 15360 19922
rect 15294 19854 15310 19888
rect 15344 19854 15360 19888
rect 15294 19820 15360 19854
rect 15294 19786 15310 19820
rect 15344 19786 15360 19820
rect 15294 19752 15360 19786
rect 15294 19718 15310 19752
rect 15344 19718 15360 19752
rect 15294 19684 15360 19718
rect 15294 19650 15310 19684
rect 15344 19650 15360 19684
rect 15294 19616 15360 19650
rect 15294 19582 15310 19616
rect 15344 19582 15360 19616
rect 15294 19548 15360 19582
rect 15294 19514 15310 19548
rect 15344 19514 15360 19548
rect 15294 19480 15360 19514
rect 15294 19446 15310 19480
rect 15344 19446 15360 19480
rect 15294 19412 15360 19446
rect 15294 19378 15310 19412
rect 15344 19378 15360 19412
rect 15294 19344 15360 19378
rect 15294 19310 15310 19344
rect 15344 19310 15360 19344
rect 15294 19276 15360 19310
rect 15294 19242 15310 19276
rect 15344 19242 15360 19276
rect 15294 19208 15360 19242
rect 15294 19174 15310 19208
rect 15344 19174 15360 19208
rect 15294 19160 15360 19174
rect 15390 20432 15456 20446
rect 15390 20398 15406 20432
rect 15440 20398 15456 20432
rect 15390 20364 15456 20398
rect 15390 20330 15406 20364
rect 15440 20330 15456 20364
rect 15390 20296 15456 20330
rect 15390 20262 15406 20296
rect 15440 20262 15456 20296
rect 15390 20228 15456 20262
rect 15390 20194 15406 20228
rect 15440 20194 15456 20228
rect 15390 20160 15456 20194
rect 15390 20126 15406 20160
rect 15440 20126 15456 20160
rect 15390 20092 15456 20126
rect 15390 20058 15406 20092
rect 15440 20058 15456 20092
rect 15390 20024 15456 20058
rect 15390 19990 15406 20024
rect 15440 19990 15456 20024
rect 15390 19956 15456 19990
rect 15390 19922 15406 19956
rect 15440 19922 15456 19956
rect 15390 19888 15456 19922
rect 15390 19854 15406 19888
rect 15440 19854 15456 19888
rect 15390 19820 15456 19854
rect 15390 19786 15406 19820
rect 15440 19786 15456 19820
rect 15390 19752 15456 19786
rect 15390 19718 15406 19752
rect 15440 19718 15456 19752
rect 15390 19684 15456 19718
rect 15390 19650 15406 19684
rect 15440 19650 15456 19684
rect 15390 19616 15456 19650
rect 15390 19582 15406 19616
rect 15440 19582 15456 19616
rect 15390 19548 15456 19582
rect 15390 19514 15406 19548
rect 15440 19514 15456 19548
rect 15390 19480 15456 19514
rect 15390 19446 15406 19480
rect 15440 19446 15456 19480
rect 15390 19412 15456 19446
rect 15390 19378 15406 19412
rect 15440 19378 15456 19412
rect 15390 19344 15456 19378
rect 15390 19310 15406 19344
rect 15440 19310 15456 19344
rect 15390 19276 15456 19310
rect 15390 19242 15406 19276
rect 15440 19242 15456 19276
rect 15390 19208 15456 19242
rect 15390 19174 15406 19208
rect 15440 19174 15456 19208
rect 15390 19160 15456 19174
rect 15486 20432 15548 20446
rect 15486 20398 15502 20432
rect 15536 20398 15548 20432
rect 15486 20364 15548 20398
rect 15486 20330 15502 20364
rect 15536 20330 15548 20364
rect 15486 20296 15548 20330
rect 15486 20262 15502 20296
rect 15536 20262 15548 20296
rect 15486 20228 15548 20262
rect 15486 20194 15502 20228
rect 15536 20194 15548 20228
rect 15486 20160 15548 20194
rect 15486 20126 15502 20160
rect 15536 20126 15548 20160
rect 15486 20092 15548 20126
rect 15486 20058 15502 20092
rect 15536 20058 15548 20092
rect 15486 20024 15548 20058
rect 15486 19990 15502 20024
rect 15536 19990 15548 20024
rect 15486 19956 15548 19990
rect 15486 19922 15502 19956
rect 15536 19922 15548 19956
rect 15486 19888 15548 19922
rect 15486 19854 15502 19888
rect 15536 19854 15548 19888
rect 15486 19820 15548 19854
rect 15486 19786 15502 19820
rect 15536 19786 15548 19820
rect 15486 19752 15548 19786
rect 15486 19718 15502 19752
rect 15536 19718 15548 19752
rect 15486 19684 15548 19718
rect 15486 19650 15502 19684
rect 15536 19650 15548 19684
rect 15486 19616 15548 19650
rect 15486 19582 15502 19616
rect 15536 19582 15548 19616
rect 15486 19548 15548 19582
rect 15486 19514 15502 19548
rect 15536 19514 15548 19548
rect 15486 19480 15548 19514
rect 15486 19446 15502 19480
rect 15536 19446 15548 19480
rect 15486 19412 15548 19446
rect 15486 19378 15502 19412
rect 15536 19378 15548 19412
rect 15486 19344 15548 19378
rect 15486 19310 15502 19344
rect 15536 19310 15548 19344
rect 15486 19276 15548 19310
rect 15486 19242 15502 19276
rect 15536 19242 15548 19276
rect 15486 19208 15548 19242
rect 15486 19174 15502 19208
rect 15536 19174 15548 19208
rect 15486 19160 15548 19174
rect 15978 19917 16040 19960
rect 15978 19883 15990 19917
rect 16024 19883 16040 19917
rect 15978 19849 16040 19883
rect 15978 19815 15990 19849
rect 16024 19815 16040 19849
rect 15978 19781 16040 19815
rect 15978 19747 15990 19781
rect 16024 19747 16040 19781
rect 15978 19713 16040 19747
rect 15978 19679 15990 19713
rect 16024 19679 16040 19713
rect 15978 19645 16040 19679
rect 15978 19611 15990 19645
rect 16024 19611 16040 19645
rect 15978 19577 16040 19611
rect 15978 19543 15990 19577
rect 16024 19543 16040 19577
rect 15978 19509 16040 19543
rect 15978 19475 15990 19509
rect 16024 19475 16040 19509
rect 15978 19441 16040 19475
rect 15978 19407 15990 19441
rect 16024 19407 16040 19441
rect 15978 19373 16040 19407
rect 15978 19339 15990 19373
rect 16024 19339 16040 19373
rect 15978 19305 16040 19339
rect 15978 19271 15990 19305
rect 16024 19271 16040 19305
rect 15978 19237 16040 19271
rect 15978 19203 15990 19237
rect 16024 19203 16040 19237
rect 15978 19160 16040 19203
rect 16070 19917 16136 19960
rect 16070 19883 16086 19917
rect 16120 19883 16136 19917
rect 16070 19849 16136 19883
rect 16070 19815 16086 19849
rect 16120 19815 16136 19849
rect 16070 19781 16136 19815
rect 16070 19747 16086 19781
rect 16120 19747 16136 19781
rect 16070 19713 16136 19747
rect 16070 19679 16086 19713
rect 16120 19679 16136 19713
rect 16070 19645 16136 19679
rect 16070 19611 16086 19645
rect 16120 19611 16136 19645
rect 16070 19577 16136 19611
rect 16070 19543 16086 19577
rect 16120 19543 16136 19577
rect 16070 19509 16136 19543
rect 16070 19475 16086 19509
rect 16120 19475 16136 19509
rect 16070 19441 16136 19475
rect 16070 19407 16086 19441
rect 16120 19407 16136 19441
rect 16070 19373 16136 19407
rect 16070 19339 16086 19373
rect 16120 19339 16136 19373
rect 16070 19305 16136 19339
rect 16070 19271 16086 19305
rect 16120 19271 16136 19305
rect 16070 19237 16136 19271
rect 16070 19203 16086 19237
rect 16120 19203 16136 19237
rect 16070 19160 16136 19203
rect 16166 19917 16232 19960
rect 16166 19883 16182 19917
rect 16216 19883 16232 19917
rect 16166 19849 16232 19883
rect 16166 19815 16182 19849
rect 16216 19815 16232 19849
rect 16166 19781 16232 19815
rect 16166 19747 16182 19781
rect 16216 19747 16232 19781
rect 16166 19713 16232 19747
rect 16166 19679 16182 19713
rect 16216 19679 16232 19713
rect 16166 19645 16232 19679
rect 16166 19611 16182 19645
rect 16216 19611 16232 19645
rect 16166 19577 16232 19611
rect 16166 19543 16182 19577
rect 16216 19543 16232 19577
rect 16166 19509 16232 19543
rect 16166 19475 16182 19509
rect 16216 19475 16232 19509
rect 16166 19441 16232 19475
rect 16166 19407 16182 19441
rect 16216 19407 16232 19441
rect 16166 19373 16232 19407
rect 16166 19339 16182 19373
rect 16216 19339 16232 19373
rect 16166 19305 16232 19339
rect 16166 19271 16182 19305
rect 16216 19271 16232 19305
rect 16166 19237 16232 19271
rect 16166 19203 16182 19237
rect 16216 19203 16232 19237
rect 16166 19160 16232 19203
rect 16262 19917 16324 19960
rect 16262 19883 16278 19917
rect 16312 19883 16324 19917
rect 16262 19849 16324 19883
rect 16262 19815 16278 19849
rect 16312 19815 16324 19849
rect 16262 19781 16324 19815
rect 16262 19747 16278 19781
rect 16312 19747 16324 19781
rect 16262 19713 16324 19747
rect 16262 19679 16278 19713
rect 16312 19679 16324 19713
rect 16262 19645 16324 19679
rect 16262 19611 16278 19645
rect 16312 19611 16324 19645
rect 16262 19577 16324 19611
rect 16262 19543 16278 19577
rect 16312 19543 16324 19577
rect 16262 19509 16324 19543
rect 16262 19475 16278 19509
rect 16312 19475 16324 19509
rect 16262 19441 16324 19475
rect 16262 19407 16278 19441
rect 16312 19407 16324 19441
rect 16262 19373 16324 19407
rect 16262 19339 16278 19373
rect 16312 19339 16324 19373
rect 16262 19305 16324 19339
rect 16262 19271 16278 19305
rect 16312 19271 16324 19305
rect 16262 19237 16324 19271
rect 16262 19203 16278 19237
rect 16312 19203 16324 19237
rect 16262 19160 16324 19203
rect 15004 18479 15062 18494
rect 15004 18445 15016 18479
rect 15050 18445 15062 18479
rect 15004 18411 15062 18445
rect 15004 18377 15016 18411
rect 15050 18377 15062 18411
rect 15004 18343 15062 18377
rect 15004 18309 15016 18343
rect 15050 18309 15062 18343
rect 15004 18275 15062 18309
rect 15004 18241 15016 18275
rect 15050 18241 15062 18275
rect 15004 18207 15062 18241
rect 15004 18173 15016 18207
rect 15050 18173 15062 18207
rect 15004 18139 15062 18173
rect 15004 18105 15016 18139
rect 15050 18105 15062 18139
rect 15004 18071 15062 18105
rect 15004 18037 15016 18071
rect 15050 18037 15062 18071
rect 15004 18003 15062 18037
rect 15004 17969 15016 18003
rect 15050 17969 15062 18003
rect 15004 17935 15062 17969
rect 15004 17901 15016 17935
rect 15050 17901 15062 17935
rect 15004 17867 15062 17901
rect 15004 17833 15016 17867
rect 15050 17833 15062 17867
rect 15004 17799 15062 17833
rect 15004 17765 15016 17799
rect 15050 17765 15062 17799
rect 15004 17731 15062 17765
rect 15004 17697 15016 17731
rect 15050 17697 15062 17731
rect 15004 17663 15062 17697
rect 15004 17629 15016 17663
rect 15050 17629 15062 17663
rect 15004 17595 15062 17629
rect 15004 17561 15016 17595
rect 15050 17561 15062 17595
rect 15004 17527 15062 17561
rect 15004 17493 15016 17527
rect 15050 17493 15062 17527
rect 15004 17459 15062 17493
rect 15004 17425 15016 17459
rect 15050 17425 15062 17459
rect 15004 17391 15062 17425
rect 15004 17357 15016 17391
rect 15050 17357 15062 17391
rect 15004 17323 15062 17357
rect 15004 17289 15016 17323
rect 15050 17289 15062 17323
rect 15004 17255 15062 17289
rect 15004 17221 15016 17255
rect 15050 17221 15062 17255
rect 15004 17187 15062 17221
rect 15004 17153 15016 17187
rect 15050 17153 15062 17187
rect 15004 17119 15062 17153
rect 15004 17085 15016 17119
rect 15050 17085 15062 17119
rect 15004 17051 15062 17085
rect 15004 17017 15016 17051
rect 15050 17017 15062 17051
rect 15004 16983 15062 17017
rect 15004 16949 15016 16983
rect 15050 16949 15062 16983
rect 15004 16934 15062 16949
rect 15092 18479 15150 18494
rect 15092 18445 15104 18479
rect 15138 18445 15150 18479
rect 15092 18411 15150 18445
rect 15092 18377 15104 18411
rect 15138 18377 15150 18411
rect 15092 18343 15150 18377
rect 15092 18309 15104 18343
rect 15138 18309 15150 18343
rect 15092 18275 15150 18309
rect 15092 18241 15104 18275
rect 15138 18241 15150 18275
rect 15092 18207 15150 18241
rect 15092 18173 15104 18207
rect 15138 18173 15150 18207
rect 15092 18139 15150 18173
rect 15092 18105 15104 18139
rect 15138 18105 15150 18139
rect 15092 18071 15150 18105
rect 15092 18037 15104 18071
rect 15138 18037 15150 18071
rect 15092 18003 15150 18037
rect 15092 17969 15104 18003
rect 15138 17969 15150 18003
rect 15092 17935 15150 17969
rect 15092 17901 15104 17935
rect 15138 17901 15150 17935
rect 15092 17867 15150 17901
rect 15092 17833 15104 17867
rect 15138 17833 15150 17867
rect 15092 17799 15150 17833
rect 15092 17765 15104 17799
rect 15138 17765 15150 17799
rect 15092 17731 15150 17765
rect 15092 17697 15104 17731
rect 15138 17697 15150 17731
rect 15092 17663 15150 17697
rect 15092 17629 15104 17663
rect 15138 17629 15150 17663
rect 15092 17595 15150 17629
rect 15092 17561 15104 17595
rect 15138 17561 15150 17595
rect 15092 17527 15150 17561
rect 15092 17493 15104 17527
rect 15138 17493 15150 17527
rect 15092 17459 15150 17493
rect 15092 17425 15104 17459
rect 15138 17425 15150 17459
rect 15092 17391 15150 17425
rect 15092 17357 15104 17391
rect 15138 17357 15150 17391
rect 15092 17323 15150 17357
rect 15092 17289 15104 17323
rect 15138 17289 15150 17323
rect 15092 17255 15150 17289
rect 15092 17221 15104 17255
rect 15138 17221 15150 17255
rect 15092 17187 15150 17221
rect 15092 17153 15104 17187
rect 15138 17153 15150 17187
rect 15092 17119 15150 17153
rect 15092 17085 15104 17119
rect 15138 17085 15150 17119
rect 15092 17051 15150 17085
rect 15092 17017 15104 17051
rect 15138 17017 15150 17051
rect 15092 16983 15150 17017
rect 15092 16949 15104 16983
rect 15138 16949 15150 16983
rect 15092 16934 15150 16949
rect 15414 18479 15472 18494
rect 15414 18445 15426 18479
rect 15460 18445 15472 18479
rect 15414 18411 15472 18445
rect 15414 18377 15426 18411
rect 15460 18377 15472 18411
rect 15414 18343 15472 18377
rect 15414 18309 15426 18343
rect 15460 18309 15472 18343
rect 15414 18275 15472 18309
rect 15414 18241 15426 18275
rect 15460 18241 15472 18275
rect 15414 18207 15472 18241
rect 15414 18173 15426 18207
rect 15460 18173 15472 18207
rect 15414 18139 15472 18173
rect 15414 18105 15426 18139
rect 15460 18105 15472 18139
rect 15414 18071 15472 18105
rect 15414 18037 15426 18071
rect 15460 18037 15472 18071
rect 15414 18003 15472 18037
rect 15414 17969 15426 18003
rect 15460 17969 15472 18003
rect 15414 17935 15472 17969
rect 15414 17901 15426 17935
rect 15460 17901 15472 17935
rect 15414 17867 15472 17901
rect 15414 17833 15426 17867
rect 15460 17833 15472 17867
rect 15414 17799 15472 17833
rect 15414 17765 15426 17799
rect 15460 17765 15472 17799
rect 15414 17731 15472 17765
rect 15414 17697 15426 17731
rect 15460 17697 15472 17731
rect 15414 17663 15472 17697
rect 15414 17629 15426 17663
rect 15460 17629 15472 17663
rect 15414 17595 15472 17629
rect 15414 17561 15426 17595
rect 15460 17561 15472 17595
rect 15414 17527 15472 17561
rect 15414 17493 15426 17527
rect 15460 17493 15472 17527
rect 15414 17459 15472 17493
rect 15414 17425 15426 17459
rect 15460 17425 15472 17459
rect 15414 17391 15472 17425
rect 15414 17357 15426 17391
rect 15460 17357 15472 17391
rect 15414 17323 15472 17357
rect 15414 17289 15426 17323
rect 15460 17289 15472 17323
rect 15414 17255 15472 17289
rect 15414 17221 15426 17255
rect 15460 17221 15472 17255
rect 15414 17187 15472 17221
rect 15414 17153 15426 17187
rect 15460 17153 15472 17187
rect 15414 17119 15472 17153
rect 15414 17085 15426 17119
rect 15460 17085 15472 17119
rect 15414 17051 15472 17085
rect 15414 17017 15426 17051
rect 15460 17017 15472 17051
rect 15414 16983 15472 17017
rect 15414 16949 15426 16983
rect 15460 16949 15472 16983
rect 15414 16934 15472 16949
rect 15502 18479 15560 18494
rect 15502 18445 15514 18479
rect 15548 18445 15560 18479
rect 15502 18411 15560 18445
rect 15502 18377 15514 18411
rect 15548 18377 15560 18411
rect 15502 18343 15560 18377
rect 15502 18309 15514 18343
rect 15548 18309 15560 18343
rect 15502 18275 15560 18309
rect 15502 18241 15514 18275
rect 15548 18241 15560 18275
rect 15502 18207 15560 18241
rect 15502 18173 15514 18207
rect 15548 18173 15560 18207
rect 15502 18139 15560 18173
rect 15502 18105 15514 18139
rect 15548 18105 15560 18139
rect 15502 18071 15560 18105
rect 15502 18037 15514 18071
rect 15548 18037 15560 18071
rect 15502 18003 15560 18037
rect 15502 17969 15514 18003
rect 15548 17969 15560 18003
rect 15502 17935 15560 17969
rect 15502 17901 15514 17935
rect 15548 17901 15560 17935
rect 15502 17867 15560 17901
rect 15502 17833 15514 17867
rect 15548 17833 15560 17867
rect 15502 17799 15560 17833
rect 15502 17765 15514 17799
rect 15548 17765 15560 17799
rect 15502 17731 15560 17765
rect 15502 17697 15514 17731
rect 15548 17697 15560 17731
rect 15502 17663 15560 17697
rect 15502 17629 15514 17663
rect 15548 17629 15560 17663
rect 15502 17595 15560 17629
rect 15502 17561 15514 17595
rect 15548 17561 15560 17595
rect 15502 17527 15560 17561
rect 15502 17493 15514 17527
rect 15548 17493 15560 17527
rect 15502 17459 15560 17493
rect 15502 17425 15514 17459
rect 15548 17425 15560 17459
rect 15502 17391 15560 17425
rect 15502 17357 15514 17391
rect 15548 17357 15560 17391
rect 15502 17323 15560 17357
rect 15502 17289 15514 17323
rect 15548 17289 15560 17323
rect 15502 17255 15560 17289
rect 15502 17221 15514 17255
rect 15548 17221 15560 17255
rect 15502 17187 15560 17221
rect 15502 17153 15514 17187
rect 15548 17153 15560 17187
rect 15502 17119 15560 17153
rect 15502 17085 15514 17119
rect 15548 17085 15560 17119
rect 15502 17051 15560 17085
rect 15502 17017 15514 17051
rect 15548 17017 15560 17051
rect 15502 16983 15560 17017
rect 15502 16949 15514 16983
rect 15548 16949 15560 16983
rect 15502 16934 15560 16949
rect 13560 15449 13618 15464
rect 13560 15415 13572 15449
rect 13606 15415 13618 15449
rect 13560 15381 13618 15415
rect 13560 15347 13572 15381
rect 13606 15347 13618 15381
rect 13560 15313 13618 15347
rect 13560 15279 13572 15313
rect 13606 15279 13618 15313
rect 13560 15245 13618 15279
rect 13560 15211 13572 15245
rect 13606 15211 13618 15245
rect 13560 15177 13618 15211
rect 13560 15143 13572 15177
rect 13606 15143 13618 15177
rect 13560 15109 13618 15143
rect 13560 15075 13572 15109
rect 13606 15075 13618 15109
rect 13560 15041 13618 15075
rect 13560 15007 13572 15041
rect 13606 15007 13618 15041
rect 13560 14973 13618 15007
rect 13560 14939 13572 14973
rect 13606 14939 13618 14973
rect 13560 14905 13618 14939
rect 13560 14871 13572 14905
rect 13606 14871 13618 14905
rect 13560 14837 13618 14871
rect 13560 14803 13572 14837
rect 13606 14803 13618 14837
rect 13560 14769 13618 14803
rect 13560 14735 13572 14769
rect 13606 14735 13618 14769
rect 13560 14701 13618 14735
rect 13560 14667 13572 14701
rect 13606 14667 13618 14701
rect 13560 14633 13618 14667
rect 13560 14599 13572 14633
rect 13606 14599 13618 14633
rect 13560 14565 13618 14599
rect 13560 14531 13572 14565
rect 13606 14531 13618 14565
rect 13560 14497 13618 14531
rect 13560 14463 13572 14497
rect 13606 14463 13618 14497
rect 13560 14429 13618 14463
rect 13560 14395 13572 14429
rect 13606 14395 13618 14429
rect 13560 14361 13618 14395
rect 13560 14327 13572 14361
rect 13606 14327 13618 14361
rect 13560 14293 13618 14327
rect 13560 14259 13572 14293
rect 13606 14259 13618 14293
rect 13560 14225 13618 14259
rect 13560 14191 13572 14225
rect 13606 14191 13618 14225
rect 13560 14157 13618 14191
rect 13560 14123 13572 14157
rect 13606 14123 13618 14157
rect 13560 14089 13618 14123
rect 13560 14055 13572 14089
rect 13606 14055 13618 14089
rect 13560 14021 13618 14055
rect 13560 13987 13572 14021
rect 13606 13987 13618 14021
rect 13560 13953 13618 13987
rect 13560 13919 13572 13953
rect 13606 13919 13618 13953
rect 13560 13904 13618 13919
rect 13648 15449 13706 15464
rect 13648 15415 13660 15449
rect 13694 15415 13706 15449
rect 13648 15381 13706 15415
rect 13648 15347 13660 15381
rect 13694 15347 13706 15381
rect 13648 15313 13706 15347
rect 13648 15279 13660 15313
rect 13694 15279 13706 15313
rect 13648 15245 13706 15279
rect 13648 15211 13660 15245
rect 13694 15211 13706 15245
rect 13648 15177 13706 15211
rect 13648 15143 13660 15177
rect 13694 15143 13706 15177
rect 13648 15109 13706 15143
rect 13648 15075 13660 15109
rect 13694 15075 13706 15109
rect 13648 15041 13706 15075
rect 13648 15007 13660 15041
rect 13694 15007 13706 15041
rect 13648 14973 13706 15007
rect 13648 14939 13660 14973
rect 13694 14939 13706 14973
rect 13648 14905 13706 14939
rect 13648 14871 13660 14905
rect 13694 14871 13706 14905
rect 13648 14837 13706 14871
rect 13648 14803 13660 14837
rect 13694 14803 13706 14837
rect 13648 14769 13706 14803
rect 13648 14735 13660 14769
rect 13694 14735 13706 14769
rect 13648 14701 13706 14735
rect 13648 14667 13660 14701
rect 13694 14667 13706 14701
rect 13648 14633 13706 14667
rect 13648 14599 13660 14633
rect 13694 14599 13706 14633
rect 13648 14565 13706 14599
rect 13648 14531 13660 14565
rect 13694 14531 13706 14565
rect 13648 14497 13706 14531
rect 13648 14463 13660 14497
rect 13694 14463 13706 14497
rect 13648 14429 13706 14463
rect 13648 14395 13660 14429
rect 13694 14395 13706 14429
rect 13648 14361 13706 14395
rect 13648 14327 13660 14361
rect 13694 14327 13706 14361
rect 13648 14293 13706 14327
rect 13648 14259 13660 14293
rect 13694 14259 13706 14293
rect 13648 14225 13706 14259
rect 13648 14191 13660 14225
rect 13694 14191 13706 14225
rect 13648 14157 13706 14191
rect 13648 14123 13660 14157
rect 13694 14123 13706 14157
rect 13648 14089 13706 14123
rect 13648 14055 13660 14089
rect 13694 14055 13706 14089
rect 13648 14021 13706 14055
rect 13648 13987 13660 14021
rect 13694 13987 13706 14021
rect 13648 13953 13706 13987
rect 13648 13919 13660 13953
rect 13694 13919 13706 13953
rect 13648 13904 13706 13919
rect 14410 15873 14472 15904
rect 14410 15839 14422 15873
rect 14456 15839 14472 15873
rect 14410 15805 14472 15839
rect 14410 15771 14422 15805
rect 14456 15771 14472 15805
rect 14410 15737 14472 15771
rect 14410 15703 14422 15737
rect 14456 15703 14472 15737
rect 14410 15669 14472 15703
rect 14410 15635 14422 15669
rect 14456 15635 14472 15669
rect 14410 15601 14472 15635
rect 14410 15567 14422 15601
rect 14456 15567 14472 15601
rect 14410 15533 14472 15567
rect 14410 15499 14422 15533
rect 14456 15499 14472 15533
rect 14410 15465 14472 15499
rect 14410 15431 14422 15465
rect 14456 15431 14472 15465
rect 14410 15397 14472 15431
rect 14410 15363 14422 15397
rect 14456 15363 14472 15397
rect 14410 15329 14472 15363
rect 14410 15295 14422 15329
rect 14456 15295 14472 15329
rect 14410 15261 14472 15295
rect 14410 15227 14422 15261
rect 14456 15227 14472 15261
rect 14410 15193 14472 15227
rect 14410 15159 14422 15193
rect 14456 15159 14472 15193
rect 14410 15125 14472 15159
rect 14410 15091 14422 15125
rect 14456 15091 14472 15125
rect 14410 15057 14472 15091
rect 14410 15023 14422 15057
rect 14456 15023 14472 15057
rect 14410 14989 14472 15023
rect 14410 14955 14422 14989
rect 14456 14955 14472 14989
rect 14410 14921 14472 14955
rect 14410 14887 14422 14921
rect 14456 14887 14472 14921
rect 14410 14853 14472 14887
rect 14410 14819 14422 14853
rect 14456 14819 14472 14853
rect 14410 14785 14472 14819
rect 14410 14751 14422 14785
rect 14456 14751 14472 14785
rect 14410 14717 14472 14751
rect 14410 14683 14422 14717
rect 14456 14683 14472 14717
rect 14410 14649 14472 14683
rect 14410 14615 14422 14649
rect 14456 14615 14472 14649
rect 14410 14581 14472 14615
rect 14410 14547 14422 14581
rect 14456 14547 14472 14581
rect 14410 14513 14472 14547
rect 14410 14479 14422 14513
rect 14456 14479 14472 14513
rect 14410 14445 14472 14479
rect 14410 14411 14422 14445
rect 14456 14411 14472 14445
rect 14410 14377 14472 14411
rect 14410 14343 14422 14377
rect 14456 14343 14472 14377
rect 14410 14309 14472 14343
rect 14410 14275 14422 14309
rect 14456 14275 14472 14309
rect 14410 14241 14472 14275
rect 14410 14207 14422 14241
rect 14456 14207 14472 14241
rect 14410 14173 14472 14207
rect 14410 14139 14422 14173
rect 14456 14139 14472 14173
rect 14410 14105 14472 14139
rect 14410 14071 14422 14105
rect 14456 14071 14472 14105
rect 14410 14037 14472 14071
rect 14410 14003 14422 14037
rect 14456 14003 14472 14037
rect 14410 13969 14472 14003
rect 14410 13935 14422 13969
rect 14456 13935 14472 13969
rect 14410 13904 14472 13935
rect 14502 15873 14568 15904
rect 14502 15839 14518 15873
rect 14552 15839 14568 15873
rect 14502 15805 14568 15839
rect 14502 15771 14518 15805
rect 14552 15771 14568 15805
rect 14502 15737 14568 15771
rect 14502 15703 14518 15737
rect 14552 15703 14568 15737
rect 14502 15669 14568 15703
rect 14502 15635 14518 15669
rect 14552 15635 14568 15669
rect 14502 15601 14568 15635
rect 14502 15567 14518 15601
rect 14552 15567 14568 15601
rect 14502 15533 14568 15567
rect 14502 15499 14518 15533
rect 14552 15499 14568 15533
rect 14502 15465 14568 15499
rect 14502 15431 14518 15465
rect 14552 15431 14568 15465
rect 14502 15397 14568 15431
rect 14502 15363 14518 15397
rect 14552 15363 14568 15397
rect 14502 15329 14568 15363
rect 14502 15295 14518 15329
rect 14552 15295 14568 15329
rect 14502 15261 14568 15295
rect 14502 15227 14518 15261
rect 14552 15227 14568 15261
rect 14502 15193 14568 15227
rect 14502 15159 14518 15193
rect 14552 15159 14568 15193
rect 14502 15125 14568 15159
rect 14502 15091 14518 15125
rect 14552 15091 14568 15125
rect 14502 15057 14568 15091
rect 14502 15023 14518 15057
rect 14552 15023 14568 15057
rect 14502 14989 14568 15023
rect 14502 14955 14518 14989
rect 14552 14955 14568 14989
rect 14502 14921 14568 14955
rect 14502 14887 14518 14921
rect 14552 14887 14568 14921
rect 14502 14853 14568 14887
rect 14502 14819 14518 14853
rect 14552 14819 14568 14853
rect 14502 14785 14568 14819
rect 14502 14751 14518 14785
rect 14552 14751 14568 14785
rect 14502 14717 14568 14751
rect 14502 14683 14518 14717
rect 14552 14683 14568 14717
rect 14502 14649 14568 14683
rect 14502 14615 14518 14649
rect 14552 14615 14568 14649
rect 14502 14581 14568 14615
rect 14502 14547 14518 14581
rect 14552 14547 14568 14581
rect 14502 14513 14568 14547
rect 14502 14479 14518 14513
rect 14552 14479 14568 14513
rect 14502 14445 14568 14479
rect 14502 14411 14518 14445
rect 14552 14411 14568 14445
rect 14502 14377 14568 14411
rect 14502 14343 14518 14377
rect 14552 14343 14568 14377
rect 14502 14309 14568 14343
rect 14502 14275 14518 14309
rect 14552 14275 14568 14309
rect 14502 14241 14568 14275
rect 14502 14207 14518 14241
rect 14552 14207 14568 14241
rect 14502 14173 14568 14207
rect 14502 14139 14518 14173
rect 14552 14139 14568 14173
rect 14502 14105 14568 14139
rect 14502 14071 14518 14105
rect 14552 14071 14568 14105
rect 14502 14037 14568 14071
rect 14502 14003 14518 14037
rect 14552 14003 14568 14037
rect 14502 13969 14568 14003
rect 14502 13935 14518 13969
rect 14552 13935 14568 13969
rect 14502 13904 14568 13935
rect 14598 15873 14664 15904
rect 14598 15839 14614 15873
rect 14648 15839 14664 15873
rect 14598 15805 14664 15839
rect 14598 15771 14614 15805
rect 14648 15771 14664 15805
rect 14598 15737 14664 15771
rect 14598 15703 14614 15737
rect 14648 15703 14664 15737
rect 14598 15669 14664 15703
rect 14598 15635 14614 15669
rect 14648 15635 14664 15669
rect 14598 15601 14664 15635
rect 14598 15567 14614 15601
rect 14648 15567 14664 15601
rect 14598 15533 14664 15567
rect 14598 15499 14614 15533
rect 14648 15499 14664 15533
rect 14598 15465 14664 15499
rect 14598 15431 14614 15465
rect 14648 15431 14664 15465
rect 14598 15397 14664 15431
rect 14598 15363 14614 15397
rect 14648 15363 14664 15397
rect 14598 15329 14664 15363
rect 14598 15295 14614 15329
rect 14648 15295 14664 15329
rect 14598 15261 14664 15295
rect 14598 15227 14614 15261
rect 14648 15227 14664 15261
rect 14598 15193 14664 15227
rect 14598 15159 14614 15193
rect 14648 15159 14664 15193
rect 14598 15125 14664 15159
rect 14598 15091 14614 15125
rect 14648 15091 14664 15125
rect 14598 15057 14664 15091
rect 14598 15023 14614 15057
rect 14648 15023 14664 15057
rect 14598 14989 14664 15023
rect 14598 14955 14614 14989
rect 14648 14955 14664 14989
rect 14598 14921 14664 14955
rect 14598 14887 14614 14921
rect 14648 14887 14664 14921
rect 14598 14853 14664 14887
rect 14598 14819 14614 14853
rect 14648 14819 14664 14853
rect 14598 14785 14664 14819
rect 14598 14751 14614 14785
rect 14648 14751 14664 14785
rect 14598 14717 14664 14751
rect 14598 14683 14614 14717
rect 14648 14683 14664 14717
rect 14598 14649 14664 14683
rect 14598 14615 14614 14649
rect 14648 14615 14664 14649
rect 14598 14581 14664 14615
rect 14598 14547 14614 14581
rect 14648 14547 14664 14581
rect 14598 14513 14664 14547
rect 14598 14479 14614 14513
rect 14648 14479 14664 14513
rect 14598 14445 14664 14479
rect 14598 14411 14614 14445
rect 14648 14411 14664 14445
rect 14598 14377 14664 14411
rect 14598 14343 14614 14377
rect 14648 14343 14664 14377
rect 14598 14309 14664 14343
rect 14598 14275 14614 14309
rect 14648 14275 14664 14309
rect 14598 14241 14664 14275
rect 14598 14207 14614 14241
rect 14648 14207 14664 14241
rect 14598 14173 14664 14207
rect 14598 14139 14614 14173
rect 14648 14139 14664 14173
rect 14598 14105 14664 14139
rect 14598 14071 14614 14105
rect 14648 14071 14664 14105
rect 14598 14037 14664 14071
rect 14598 14003 14614 14037
rect 14648 14003 14664 14037
rect 14598 13969 14664 14003
rect 14598 13935 14614 13969
rect 14648 13935 14664 13969
rect 14598 13904 14664 13935
rect 14694 15873 14760 15904
rect 14694 15839 14710 15873
rect 14744 15839 14760 15873
rect 14694 15805 14760 15839
rect 14694 15771 14710 15805
rect 14744 15771 14760 15805
rect 14694 15737 14760 15771
rect 14694 15703 14710 15737
rect 14744 15703 14760 15737
rect 14694 15669 14760 15703
rect 14694 15635 14710 15669
rect 14744 15635 14760 15669
rect 14694 15601 14760 15635
rect 14694 15567 14710 15601
rect 14744 15567 14760 15601
rect 14694 15533 14760 15567
rect 14694 15499 14710 15533
rect 14744 15499 14760 15533
rect 14694 15465 14760 15499
rect 14694 15431 14710 15465
rect 14744 15431 14760 15465
rect 14694 15397 14760 15431
rect 14694 15363 14710 15397
rect 14744 15363 14760 15397
rect 14694 15329 14760 15363
rect 14694 15295 14710 15329
rect 14744 15295 14760 15329
rect 14694 15261 14760 15295
rect 14694 15227 14710 15261
rect 14744 15227 14760 15261
rect 14694 15193 14760 15227
rect 14694 15159 14710 15193
rect 14744 15159 14760 15193
rect 14694 15125 14760 15159
rect 14694 15091 14710 15125
rect 14744 15091 14760 15125
rect 14694 15057 14760 15091
rect 14694 15023 14710 15057
rect 14744 15023 14760 15057
rect 14694 14989 14760 15023
rect 14694 14955 14710 14989
rect 14744 14955 14760 14989
rect 14694 14921 14760 14955
rect 14694 14887 14710 14921
rect 14744 14887 14760 14921
rect 14694 14853 14760 14887
rect 14694 14819 14710 14853
rect 14744 14819 14760 14853
rect 14694 14785 14760 14819
rect 14694 14751 14710 14785
rect 14744 14751 14760 14785
rect 14694 14717 14760 14751
rect 14694 14683 14710 14717
rect 14744 14683 14760 14717
rect 14694 14649 14760 14683
rect 14694 14615 14710 14649
rect 14744 14615 14760 14649
rect 14694 14581 14760 14615
rect 14694 14547 14710 14581
rect 14744 14547 14760 14581
rect 14694 14513 14760 14547
rect 14694 14479 14710 14513
rect 14744 14479 14760 14513
rect 14694 14445 14760 14479
rect 14694 14411 14710 14445
rect 14744 14411 14760 14445
rect 14694 14377 14760 14411
rect 14694 14343 14710 14377
rect 14744 14343 14760 14377
rect 14694 14309 14760 14343
rect 14694 14275 14710 14309
rect 14744 14275 14760 14309
rect 14694 14241 14760 14275
rect 14694 14207 14710 14241
rect 14744 14207 14760 14241
rect 14694 14173 14760 14207
rect 14694 14139 14710 14173
rect 14744 14139 14760 14173
rect 14694 14105 14760 14139
rect 14694 14071 14710 14105
rect 14744 14071 14760 14105
rect 14694 14037 14760 14071
rect 14694 14003 14710 14037
rect 14744 14003 14760 14037
rect 14694 13969 14760 14003
rect 14694 13935 14710 13969
rect 14744 13935 14760 13969
rect 14694 13904 14760 13935
rect 14790 15873 14856 15904
rect 14790 15839 14806 15873
rect 14840 15839 14856 15873
rect 14790 15805 14856 15839
rect 14790 15771 14806 15805
rect 14840 15771 14856 15805
rect 14790 15737 14856 15771
rect 14790 15703 14806 15737
rect 14840 15703 14856 15737
rect 14790 15669 14856 15703
rect 14790 15635 14806 15669
rect 14840 15635 14856 15669
rect 14790 15601 14856 15635
rect 14790 15567 14806 15601
rect 14840 15567 14856 15601
rect 14790 15533 14856 15567
rect 14790 15499 14806 15533
rect 14840 15499 14856 15533
rect 14790 15465 14856 15499
rect 14790 15431 14806 15465
rect 14840 15431 14856 15465
rect 14790 15397 14856 15431
rect 14790 15363 14806 15397
rect 14840 15363 14856 15397
rect 14790 15329 14856 15363
rect 14790 15295 14806 15329
rect 14840 15295 14856 15329
rect 14790 15261 14856 15295
rect 14790 15227 14806 15261
rect 14840 15227 14856 15261
rect 14790 15193 14856 15227
rect 14790 15159 14806 15193
rect 14840 15159 14856 15193
rect 14790 15125 14856 15159
rect 14790 15091 14806 15125
rect 14840 15091 14856 15125
rect 14790 15057 14856 15091
rect 14790 15023 14806 15057
rect 14840 15023 14856 15057
rect 14790 14989 14856 15023
rect 14790 14955 14806 14989
rect 14840 14955 14856 14989
rect 14790 14921 14856 14955
rect 14790 14887 14806 14921
rect 14840 14887 14856 14921
rect 14790 14853 14856 14887
rect 14790 14819 14806 14853
rect 14840 14819 14856 14853
rect 14790 14785 14856 14819
rect 14790 14751 14806 14785
rect 14840 14751 14856 14785
rect 14790 14717 14856 14751
rect 14790 14683 14806 14717
rect 14840 14683 14856 14717
rect 14790 14649 14856 14683
rect 14790 14615 14806 14649
rect 14840 14615 14856 14649
rect 14790 14581 14856 14615
rect 14790 14547 14806 14581
rect 14840 14547 14856 14581
rect 14790 14513 14856 14547
rect 14790 14479 14806 14513
rect 14840 14479 14856 14513
rect 14790 14445 14856 14479
rect 14790 14411 14806 14445
rect 14840 14411 14856 14445
rect 14790 14377 14856 14411
rect 14790 14343 14806 14377
rect 14840 14343 14856 14377
rect 14790 14309 14856 14343
rect 14790 14275 14806 14309
rect 14840 14275 14856 14309
rect 14790 14241 14856 14275
rect 14790 14207 14806 14241
rect 14840 14207 14856 14241
rect 14790 14173 14856 14207
rect 14790 14139 14806 14173
rect 14840 14139 14856 14173
rect 14790 14105 14856 14139
rect 14790 14071 14806 14105
rect 14840 14071 14856 14105
rect 14790 14037 14856 14071
rect 14790 14003 14806 14037
rect 14840 14003 14856 14037
rect 14790 13969 14856 14003
rect 14790 13935 14806 13969
rect 14840 13935 14856 13969
rect 14790 13904 14856 13935
rect 14886 15873 14952 15904
rect 14886 15839 14902 15873
rect 14936 15839 14952 15873
rect 14886 15805 14952 15839
rect 14886 15771 14902 15805
rect 14936 15771 14952 15805
rect 14886 15737 14952 15771
rect 14886 15703 14902 15737
rect 14936 15703 14952 15737
rect 14886 15669 14952 15703
rect 14886 15635 14902 15669
rect 14936 15635 14952 15669
rect 14886 15601 14952 15635
rect 14886 15567 14902 15601
rect 14936 15567 14952 15601
rect 14886 15533 14952 15567
rect 14886 15499 14902 15533
rect 14936 15499 14952 15533
rect 14886 15465 14952 15499
rect 14886 15431 14902 15465
rect 14936 15431 14952 15465
rect 14886 15397 14952 15431
rect 14886 15363 14902 15397
rect 14936 15363 14952 15397
rect 14886 15329 14952 15363
rect 14886 15295 14902 15329
rect 14936 15295 14952 15329
rect 14886 15261 14952 15295
rect 14886 15227 14902 15261
rect 14936 15227 14952 15261
rect 14886 15193 14952 15227
rect 14886 15159 14902 15193
rect 14936 15159 14952 15193
rect 14886 15125 14952 15159
rect 14886 15091 14902 15125
rect 14936 15091 14952 15125
rect 14886 15057 14952 15091
rect 14886 15023 14902 15057
rect 14936 15023 14952 15057
rect 14886 14989 14952 15023
rect 14886 14955 14902 14989
rect 14936 14955 14952 14989
rect 14886 14921 14952 14955
rect 14886 14887 14902 14921
rect 14936 14887 14952 14921
rect 14886 14853 14952 14887
rect 14886 14819 14902 14853
rect 14936 14819 14952 14853
rect 14886 14785 14952 14819
rect 14886 14751 14902 14785
rect 14936 14751 14952 14785
rect 14886 14717 14952 14751
rect 14886 14683 14902 14717
rect 14936 14683 14952 14717
rect 14886 14649 14952 14683
rect 14886 14615 14902 14649
rect 14936 14615 14952 14649
rect 14886 14581 14952 14615
rect 14886 14547 14902 14581
rect 14936 14547 14952 14581
rect 14886 14513 14952 14547
rect 14886 14479 14902 14513
rect 14936 14479 14952 14513
rect 14886 14445 14952 14479
rect 14886 14411 14902 14445
rect 14936 14411 14952 14445
rect 14886 14377 14952 14411
rect 14886 14343 14902 14377
rect 14936 14343 14952 14377
rect 14886 14309 14952 14343
rect 14886 14275 14902 14309
rect 14936 14275 14952 14309
rect 14886 14241 14952 14275
rect 14886 14207 14902 14241
rect 14936 14207 14952 14241
rect 14886 14173 14952 14207
rect 14886 14139 14902 14173
rect 14936 14139 14952 14173
rect 14886 14105 14952 14139
rect 14886 14071 14902 14105
rect 14936 14071 14952 14105
rect 14886 14037 14952 14071
rect 14886 14003 14902 14037
rect 14936 14003 14952 14037
rect 14886 13969 14952 14003
rect 14886 13935 14902 13969
rect 14936 13935 14952 13969
rect 14886 13904 14952 13935
rect 14982 15873 15048 15904
rect 14982 15839 14998 15873
rect 15032 15839 15048 15873
rect 14982 15805 15048 15839
rect 14982 15771 14998 15805
rect 15032 15771 15048 15805
rect 14982 15737 15048 15771
rect 14982 15703 14998 15737
rect 15032 15703 15048 15737
rect 14982 15669 15048 15703
rect 14982 15635 14998 15669
rect 15032 15635 15048 15669
rect 14982 15601 15048 15635
rect 14982 15567 14998 15601
rect 15032 15567 15048 15601
rect 14982 15533 15048 15567
rect 14982 15499 14998 15533
rect 15032 15499 15048 15533
rect 14982 15465 15048 15499
rect 14982 15431 14998 15465
rect 15032 15431 15048 15465
rect 14982 15397 15048 15431
rect 14982 15363 14998 15397
rect 15032 15363 15048 15397
rect 14982 15329 15048 15363
rect 14982 15295 14998 15329
rect 15032 15295 15048 15329
rect 14982 15261 15048 15295
rect 14982 15227 14998 15261
rect 15032 15227 15048 15261
rect 14982 15193 15048 15227
rect 14982 15159 14998 15193
rect 15032 15159 15048 15193
rect 14982 15125 15048 15159
rect 14982 15091 14998 15125
rect 15032 15091 15048 15125
rect 14982 15057 15048 15091
rect 14982 15023 14998 15057
rect 15032 15023 15048 15057
rect 14982 14989 15048 15023
rect 14982 14955 14998 14989
rect 15032 14955 15048 14989
rect 14982 14921 15048 14955
rect 14982 14887 14998 14921
rect 15032 14887 15048 14921
rect 14982 14853 15048 14887
rect 14982 14819 14998 14853
rect 15032 14819 15048 14853
rect 14982 14785 15048 14819
rect 14982 14751 14998 14785
rect 15032 14751 15048 14785
rect 14982 14717 15048 14751
rect 14982 14683 14998 14717
rect 15032 14683 15048 14717
rect 14982 14649 15048 14683
rect 14982 14615 14998 14649
rect 15032 14615 15048 14649
rect 14982 14581 15048 14615
rect 14982 14547 14998 14581
rect 15032 14547 15048 14581
rect 14982 14513 15048 14547
rect 14982 14479 14998 14513
rect 15032 14479 15048 14513
rect 14982 14445 15048 14479
rect 14982 14411 14998 14445
rect 15032 14411 15048 14445
rect 14982 14377 15048 14411
rect 14982 14343 14998 14377
rect 15032 14343 15048 14377
rect 14982 14309 15048 14343
rect 14982 14275 14998 14309
rect 15032 14275 15048 14309
rect 14982 14241 15048 14275
rect 14982 14207 14998 14241
rect 15032 14207 15048 14241
rect 14982 14173 15048 14207
rect 14982 14139 14998 14173
rect 15032 14139 15048 14173
rect 14982 14105 15048 14139
rect 14982 14071 14998 14105
rect 15032 14071 15048 14105
rect 14982 14037 15048 14071
rect 14982 14003 14998 14037
rect 15032 14003 15048 14037
rect 14982 13969 15048 14003
rect 14982 13935 14998 13969
rect 15032 13935 15048 13969
rect 14982 13904 15048 13935
rect 15078 15873 15144 15904
rect 15078 15839 15094 15873
rect 15128 15839 15144 15873
rect 15078 15805 15144 15839
rect 15078 15771 15094 15805
rect 15128 15771 15144 15805
rect 15078 15737 15144 15771
rect 15078 15703 15094 15737
rect 15128 15703 15144 15737
rect 15078 15669 15144 15703
rect 15078 15635 15094 15669
rect 15128 15635 15144 15669
rect 15078 15601 15144 15635
rect 15078 15567 15094 15601
rect 15128 15567 15144 15601
rect 15078 15533 15144 15567
rect 15078 15499 15094 15533
rect 15128 15499 15144 15533
rect 15078 15465 15144 15499
rect 15078 15431 15094 15465
rect 15128 15431 15144 15465
rect 15078 15397 15144 15431
rect 15078 15363 15094 15397
rect 15128 15363 15144 15397
rect 15078 15329 15144 15363
rect 15078 15295 15094 15329
rect 15128 15295 15144 15329
rect 15078 15261 15144 15295
rect 15078 15227 15094 15261
rect 15128 15227 15144 15261
rect 15078 15193 15144 15227
rect 15078 15159 15094 15193
rect 15128 15159 15144 15193
rect 15078 15125 15144 15159
rect 15078 15091 15094 15125
rect 15128 15091 15144 15125
rect 15078 15057 15144 15091
rect 15078 15023 15094 15057
rect 15128 15023 15144 15057
rect 15078 14989 15144 15023
rect 15078 14955 15094 14989
rect 15128 14955 15144 14989
rect 15078 14921 15144 14955
rect 15078 14887 15094 14921
rect 15128 14887 15144 14921
rect 15078 14853 15144 14887
rect 15078 14819 15094 14853
rect 15128 14819 15144 14853
rect 15078 14785 15144 14819
rect 15078 14751 15094 14785
rect 15128 14751 15144 14785
rect 15078 14717 15144 14751
rect 15078 14683 15094 14717
rect 15128 14683 15144 14717
rect 15078 14649 15144 14683
rect 15078 14615 15094 14649
rect 15128 14615 15144 14649
rect 15078 14581 15144 14615
rect 15078 14547 15094 14581
rect 15128 14547 15144 14581
rect 15078 14513 15144 14547
rect 15078 14479 15094 14513
rect 15128 14479 15144 14513
rect 15078 14445 15144 14479
rect 15078 14411 15094 14445
rect 15128 14411 15144 14445
rect 15078 14377 15144 14411
rect 15078 14343 15094 14377
rect 15128 14343 15144 14377
rect 15078 14309 15144 14343
rect 15078 14275 15094 14309
rect 15128 14275 15144 14309
rect 15078 14241 15144 14275
rect 15078 14207 15094 14241
rect 15128 14207 15144 14241
rect 15078 14173 15144 14207
rect 15078 14139 15094 14173
rect 15128 14139 15144 14173
rect 15078 14105 15144 14139
rect 15078 14071 15094 14105
rect 15128 14071 15144 14105
rect 15078 14037 15144 14071
rect 15078 14003 15094 14037
rect 15128 14003 15144 14037
rect 15078 13969 15144 14003
rect 15078 13935 15094 13969
rect 15128 13935 15144 13969
rect 15078 13904 15144 13935
rect 15174 15873 15236 15904
rect 15174 15839 15190 15873
rect 15224 15839 15236 15873
rect 15174 15805 15236 15839
rect 15174 15771 15190 15805
rect 15224 15771 15236 15805
rect 15174 15737 15236 15771
rect 15174 15703 15190 15737
rect 15224 15703 15236 15737
rect 15174 15669 15236 15703
rect 15174 15635 15190 15669
rect 15224 15635 15236 15669
rect 15174 15601 15236 15635
rect 15174 15567 15190 15601
rect 15224 15567 15236 15601
rect 15174 15533 15236 15567
rect 15174 15499 15190 15533
rect 15224 15499 15236 15533
rect 15174 15465 15236 15499
rect 15174 15431 15190 15465
rect 15224 15431 15236 15465
rect 15174 15397 15236 15431
rect 15174 15363 15190 15397
rect 15224 15363 15236 15397
rect 15174 15329 15236 15363
rect 15174 15295 15190 15329
rect 15224 15295 15236 15329
rect 15174 15261 15236 15295
rect 15174 15227 15190 15261
rect 15224 15227 15236 15261
rect 15174 15193 15236 15227
rect 15174 15159 15190 15193
rect 15224 15159 15236 15193
rect 15174 15125 15236 15159
rect 15174 15091 15190 15125
rect 15224 15091 15236 15125
rect 15174 15057 15236 15091
rect 15174 15023 15190 15057
rect 15224 15023 15236 15057
rect 15174 14989 15236 15023
rect 15174 14955 15190 14989
rect 15224 14955 15236 14989
rect 15174 14921 15236 14955
rect 15174 14887 15190 14921
rect 15224 14887 15236 14921
rect 15174 14853 15236 14887
rect 15174 14819 15190 14853
rect 15224 14819 15236 14853
rect 15174 14785 15236 14819
rect 15174 14751 15190 14785
rect 15224 14751 15236 14785
rect 15174 14717 15236 14751
rect 15174 14683 15190 14717
rect 15224 14683 15236 14717
rect 15174 14649 15236 14683
rect 15174 14615 15190 14649
rect 15224 14615 15236 14649
rect 15174 14581 15236 14615
rect 15174 14547 15190 14581
rect 15224 14547 15236 14581
rect 15174 14513 15236 14547
rect 15174 14479 15190 14513
rect 15224 14479 15236 14513
rect 15174 14445 15236 14479
rect 15174 14411 15190 14445
rect 15224 14411 15236 14445
rect 15174 14377 15236 14411
rect 15174 14343 15190 14377
rect 15224 14343 15236 14377
rect 15174 14309 15236 14343
rect 15174 14275 15190 14309
rect 15224 14275 15236 14309
rect 15174 14241 15236 14275
rect 15174 14207 15190 14241
rect 15224 14207 15236 14241
rect 15174 14173 15236 14207
rect 15174 14139 15190 14173
rect 15224 14139 15236 14173
rect 15174 14105 15236 14139
rect 15174 14071 15190 14105
rect 15224 14071 15236 14105
rect 15174 14037 15236 14071
rect 15174 14003 15190 14037
rect 15224 14003 15236 14037
rect 15174 13969 15236 14003
rect 15174 13935 15190 13969
rect 15224 13935 15236 13969
rect 15174 13904 15236 13935
rect 13422 13039 13480 13070
rect 13422 13005 13434 13039
rect 13468 13005 13480 13039
rect 13422 12971 13480 13005
rect 13422 12937 13434 12971
rect 13468 12937 13480 12971
rect 13422 12903 13480 12937
rect 13422 12869 13434 12903
rect 13468 12869 13480 12903
rect 13422 12835 13480 12869
rect 13422 12801 13434 12835
rect 13468 12801 13480 12835
rect 13422 12767 13480 12801
rect 13422 12733 13434 12767
rect 13468 12733 13480 12767
rect 13422 12699 13480 12733
rect 13422 12665 13434 12699
rect 13468 12665 13480 12699
rect 13422 12631 13480 12665
rect 13422 12597 13434 12631
rect 13468 12597 13480 12631
rect 13422 12563 13480 12597
rect 13422 12529 13434 12563
rect 13468 12529 13480 12563
rect 13422 12495 13480 12529
rect 13422 12461 13434 12495
rect 13468 12461 13480 12495
rect 13422 12427 13480 12461
rect 13422 12393 13434 12427
rect 13468 12393 13480 12427
rect 13422 12359 13480 12393
rect 13422 12325 13434 12359
rect 13468 12325 13480 12359
rect 13422 12291 13480 12325
rect 13422 12257 13434 12291
rect 13468 12257 13480 12291
rect 13422 12223 13480 12257
rect 13422 12189 13434 12223
rect 13468 12189 13480 12223
rect 13422 12155 13480 12189
rect 13422 12121 13434 12155
rect 13468 12121 13480 12155
rect 13422 12087 13480 12121
rect 13422 12053 13434 12087
rect 13468 12053 13480 12087
rect 13422 12019 13480 12053
rect 13422 11985 13434 12019
rect 13468 11985 13480 12019
rect 13422 11951 13480 11985
rect 13422 11917 13434 11951
rect 13468 11917 13480 11951
rect 13422 11883 13480 11917
rect 13422 11849 13434 11883
rect 13468 11849 13480 11883
rect 13422 11815 13480 11849
rect 13422 11781 13434 11815
rect 13468 11781 13480 11815
rect 13422 11747 13480 11781
rect 13422 11713 13434 11747
rect 13468 11713 13480 11747
rect 13422 11679 13480 11713
rect 13422 11645 13434 11679
rect 13468 11645 13480 11679
rect 13422 11611 13480 11645
rect 13422 11577 13434 11611
rect 13468 11577 13480 11611
rect 13422 11543 13480 11577
rect 13422 11509 13434 11543
rect 13468 11509 13480 11543
rect 13422 11475 13480 11509
rect 13422 11441 13434 11475
rect 13468 11441 13480 11475
rect 13422 11407 13480 11441
rect 13422 11373 13434 11407
rect 13468 11373 13480 11407
rect 13422 11339 13480 11373
rect 13422 11305 13434 11339
rect 13468 11305 13480 11339
rect 13422 11271 13480 11305
rect 13422 11237 13434 11271
rect 13468 11237 13480 11271
rect 13422 11203 13480 11237
rect 13422 11169 13434 11203
rect 13468 11169 13480 11203
rect 13422 11135 13480 11169
rect 13422 11101 13434 11135
rect 13468 11101 13480 11135
rect 13422 11070 13480 11101
rect 13510 13039 13568 13070
rect 13510 13005 13522 13039
rect 13556 13005 13568 13039
rect 13510 12971 13568 13005
rect 13510 12937 13522 12971
rect 13556 12937 13568 12971
rect 13510 12903 13568 12937
rect 13510 12869 13522 12903
rect 13556 12869 13568 12903
rect 13510 12835 13568 12869
rect 13510 12801 13522 12835
rect 13556 12801 13568 12835
rect 13510 12767 13568 12801
rect 13510 12733 13522 12767
rect 13556 12733 13568 12767
rect 13510 12699 13568 12733
rect 13510 12665 13522 12699
rect 13556 12665 13568 12699
rect 13510 12631 13568 12665
rect 13510 12597 13522 12631
rect 13556 12597 13568 12631
rect 13510 12563 13568 12597
rect 13510 12529 13522 12563
rect 13556 12529 13568 12563
rect 13510 12495 13568 12529
rect 13510 12461 13522 12495
rect 13556 12461 13568 12495
rect 13510 12427 13568 12461
rect 13510 12393 13522 12427
rect 13556 12393 13568 12427
rect 13510 12359 13568 12393
rect 13510 12325 13522 12359
rect 13556 12325 13568 12359
rect 13510 12291 13568 12325
rect 13510 12257 13522 12291
rect 13556 12257 13568 12291
rect 13510 12223 13568 12257
rect 13510 12189 13522 12223
rect 13556 12189 13568 12223
rect 13510 12155 13568 12189
rect 13510 12121 13522 12155
rect 13556 12121 13568 12155
rect 13510 12087 13568 12121
rect 13510 12053 13522 12087
rect 13556 12053 13568 12087
rect 13510 12019 13568 12053
rect 13510 11985 13522 12019
rect 13556 11985 13568 12019
rect 13510 11951 13568 11985
rect 13510 11917 13522 11951
rect 13556 11917 13568 11951
rect 13510 11883 13568 11917
rect 13510 11849 13522 11883
rect 13556 11849 13568 11883
rect 13510 11815 13568 11849
rect 13510 11781 13522 11815
rect 13556 11781 13568 11815
rect 13510 11747 13568 11781
rect 13510 11713 13522 11747
rect 13556 11713 13568 11747
rect 13510 11679 13568 11713
rect 13510 11645 13522 11679
rect 13556 11645 13568 11679
rect 13510 11611 13568 11645
rect 13510 11577 13522 11611
rect 13556 11577 13568 11611
rect 13510 11543 13568 11577
rect 13510 11509 13522 11543
rect 13556 11509 13568 11543
rect 13510 11475 13568 11509
rect 13510 11441 13522 11475
rect 13556 11441 13568 11475
rect 13510 11407 13568 11441
rect 13510 11373 13522 11407
rect 13556 11373 13568 11407
rect 13510 11339 13568 11373
rect 13510 11305 13522 11339
rect 13556 11305 13568 11339
rect 13510 11271 13568 11305
rect 13510 11237 13522 11271
rect 13556 11237 13568 11271
rect 13510 11203 13568 11237
rect 13510 11169 13522 11203
rect 13556 11169 13568 11203
rect 13510 11135 13568 11169
rect 13510 11101 13522 11135
rect 13556 11101 13568 11135
rect 13510 11070 13568 11101
rect 13598 13039 13656 13070
rect 13598 13005 13610 13039
rect 13644 13005 13656 13039
rect 13598 12971 13656 13005
rect 13598 12937 13610 12971
rect 13644 12937 13656 12971
rect 13598 12903 13656 12937
rect 13598 12869 13610 12903
rect 13644 12869 13656 12903
rect 13598 12835 13656 12869
rect 13598 12801 13610 12835
rect 13644 12801 13656 12835
rect 13598 12767 13656 12801
rect 13598 12733 13610 12767
rect 13644 12733 13656 12767
rect 13598 12699 13656 12733
rect 13598 12665 13610 12699
rect 13644 12665 13656 12699
rect 13598 12631 13656 12665
rect 13598 12597 13610 12631
rect 13644 12597 13656 12631
rect 13598 12563 13656 12597
rect 13598 12529 13610 12563
rect 13644 12529 13656 12563
rect 13598 12495 13656 12529
rect 13598 12461 13610 12495
rect 13644 12461 13656 12495
rect 13598 12427 13656 12461
rect 13598 12393 13610 12427
rect 13644 12393 13656 12427
rect 13598 12359 13656 12393
rect 13598 12325 13610 12359
rect 13644 12325 13656 12359
rect 13598 12291 13656 12325
rect 13598 12257 13610 12291
rect 13644 12257 13656 12291
rect 13598 12223 13656 12257
rect 13598 12189 13610 12223
rect 13644 12189 13656 12223
rect 13598 12155 13656 12189
rect 13598 12121 13610 12155
rect 13644 12121 13656 12155
rect 13598 12087 13656 12121
rect 13598 12053 13610 12087
rect 13644 12053 13656 12087
rect 13598 12019 13656 12053
rect 13598 11985 13610 12019
rect 13644 11985 13656 12019
rect 13598 11951 13656 11985
rect 13598 11917 13610 11951
rect 13644 11917 13656 11951
rect 13598 11883 13656 11917
rect 13598 11849 13610 11883
rect 13644 11849 13656 11883
rect 13598 11815 13656 11849
rect 13598 11781 13610 11815
rect 13644 11781 13656 11815
rect 13598 11747 13656 11781
rect 13598 11713 13610 11747
rect 13644 11713 13656 11747
rect 13598 11679 13656 11713
rect 13598 11645 13610 11679
rect 13644 11645 13656 11679
rect 13598 11611 13656 11645
rect 13598 11577 13610 11611
rect 13644 11577 13656 11611
rect 13598 11543 13656 11577
rect 13598 11509 13610 11543
rect 13644 11509 13656 11543
rect 13598 11475 13656 11509
rect 13598 11441 13610 11475
rect 13644 11441 13656 11475
rect 13598 11407 13656 11441
rect 13598 11373 13610 11407
rect 13644 11373 13656 11407
rect 13598 11339 13656 11373
rect 13598 11305 13610 11339
rect 13644 11305 13656 11339
rect 13598 11271 13656 11305
rect 13598 11237 13610 11271
rect 13644 11237 13656 11271
rect 13598 11203 13656 11237
rect 13598 11169 13610 11203
rect 13644 11169 13656 11203
rect 13598 11135 13656 11169
rect 13598 11101 13610 11135
rect 13644 11101 13656 11135
rect 13598 11070 13656 11101
rect 13686 13039 13744 13070
rect 13686 13005 13698 13039
rect 13732 13005 13744 13039
rect 13686 12971 13744 13005
rect 13686 12937 13698 12971
rect 13732 12937 13744 12971
rect 13686 12903 13744 12937
rect 13686 12869 13698 12903
rect 13732 12869 13744 12903
rect 13686 12835 13744 12869
rect 13686 12801 13698 12835
rect 13732 12801 13744 12835
rect 13686 12767 13744 12801
rect 13686 12733 13698 12767
rect 13732 12733 13744 12767
rect 13686 12699 13744 12733
rect 13686 12665 13698 12699
rect 13732 12665 13744 12699
rect 13686 12631 13744 12665
rect 13686 12597 13698 12631
rect 13732 12597 13744 12631
rect 13686 12563 13744 12597
rect 13686 12529 13698 12563
rect 13732 12529 13744 12563
rect 13686 12495 13744 12529
rect 13686 12461 13698 12495
rect 13732 12461 13744 12495
rect 13686 12427 13744 12461
rect 13686 12393 13698 12427
rect 13732 12393 13744 12427
rect 13686 12359 13744 12393
rect 13686 12325 13698 12359
rect 13732 12325 13744 12359
rect 13686 12291 13744 12325
rect 13686 12257 13698 12291
rect 13732 12257 13744 12291
rect 13686 12223 13744 12257
rect 13686 12189 13698 12223
rect 13732 12189 13744 12223
rect 13686 12155 13744 12189
rect 13686 12121 13698 12155
rect 13732 12121 13744 12155
rect 13686 12087 13744 12121
rect 13686 12053 13698 12087
rect 13732 12053 13744 12087
rect 13686 12019 13744 12053
rect 13686 11985 13698 12019
rect 13732 11985 13744 12019
rect 13686 11951 13744 11985
rect 13686 11917 13698 11951
rect 13732 11917 13744 11951
rect 13686 11883 13744 11917
rect 13686 11849 13698 11883
rect 13732 11849 13744 11883
rect 13686 11815 13744 11849
rect 13686 11781 13698 11815
rect 13732 11781 13744 11815
rect 13686 11747 13744 11781
rect 13686 11713 13698 11747
rect 13732 11713 13744 11747
rect 13686 11679 13744 11713
rect 13686 11645 13698 11679
rect 13732 11645 13744 11679
rect 13686 11611 13744 11645
rect 13686 11577 13698 11611
rect 13732 11577 13744 11611
rect 13686 11543 13744 11577
rect 13686 11509 13698 11543
rect 13732 11509 13744 11543
rect 13686 11475 13744 11509
rect 13686 11441 13698 11475
rect 13732 11441 13744 11475
rect 13686 11407 13744 11441
rect 13686 11373 13698 11407
rect 13732 11373 13744 11407
rect 13686 11339 13744 11373
rect 13686 11305 13698 11339
rect 13732 11305 13744 11339
rect 13686 11271 13744 11305
rect 13686 11237 13698 11271
rect 13732 11237 13744 11271
rect 13686 11203 13744 11237
rect 13686 11169 13698 11203
rect 13732 11169 13744 11203
rect 13686 11135 13744 11169
rect 13686 11101 13698 11135
rect 13732 11101 13744 11135
rect 13686 11070 13744 11101
rect 13774 13039 13832 13070
rect 13774 13005 13786 13039
rect 13820 13005 13832 13039
rect 13774 12971 13832 13005
rect 13774 12937 13786 12971
rect 13820 12937 13832 12971
rect 13774 12903 13832 12937
rect 13774 12869 13786 12903
rect 13820 12869 13832 12903
rect 13774 12835 13832 12869
rect 13774 12801 13786 12835
rect 13820 12801 13832 12835
rect 13774 12767 13832 12801
rect 13774 12733 13786 12767
rect 13820 12733 13832 12767
rect 13774 12699 13832 12733
rect 13774 12665 13786 12699
rect 13820 12665 13832 12699
rect 13774 12631 13832 12665
rect 13774 12597 13786 12631
rect 13820 12597 13832 12631
rect 13774 12563 13832 12597
rect 13774 12529 13786 12563
rect 13820 12529 13832 12563
rect 13774 12495 13832 12529
rect 13774 12461 13786 12495
rect 13820 12461 13832 12495
rect 13774 12427 13832 12461
rect 13774 12393 13786 12427
rect 13820 12393 13832 12427
rect 13774 12359 13832 12393
rect 13774 12325 13786 12359
rect 13820 12325 13832 12359
rect 13774 12291 13832 12325
rect 13774 12257 13786 12291
rect 13820 12257 13832 12291
rect 13774 12223 13832 12257
rect 13774 12189 13786 12223
rect 13820 12189 13832 12223
rect 13774 12155 13832 12189
rect 13774 12121 13786 12155
rect 13820 12121 13832 12155
rect 13774 12087 13832 12121
rect 13774 12053 13786 12087
rect 13820 12053 13832 12087
rect 13774 12019 13832 12053
rect 13774 11985 13786 12019
rect 13820 11985 13832 12019
rect 13774 11951 13832 11985
rect 13774 11917 13786 11951
rect 13820 11917 13832 11951
rect 13774 11883 13832 11917
rect 13774 11849 13786 11883
rect 13820 11849 13832 11883
rect 13774 11815 13832 11849
rect 13774 11781 13786 11815
rect 13820 11781 13832 11815
rect 13774 11747 13832 11781
rect 13774 11713 13786 11747
rect 13820 11713 13832 11747
rect 13774 11679 13832 11713
rect 13774 11645 13786 11679
rect 13820 11645 13832 11679
rect 13774 11611 13832 11645
rect 13774 11577 13786 11611
rect 13820 11577 13832 11611
rect 13774 11543 13832 11577
rect 13774 11509 13786 11543
rect 13820 11509 13832 11543
rect 13774 11475 13832 11509
rect 13774 11441 13786 11475
rect 13820 11441 13832 11475
rect 13774 11407 13832 11441
rect 13774 11373 13786 11407
rect 13820 11373 13832 11407
rect 13774 11339 13832 11373
rect 13774 11305 13786 11339
rect 13820 11305 13832 11339
rect 13774 11271 13832 11305
rect 13774 11237 13786 11271
rect 13820 11237 13832 11271
rect 13774 11203 13832 11237
rect 13774 11169 13786 11203
rect 13820 11169 13832 11203
rect 13774 11135 13832 11169
rect 13774 11101 13786 11135
rect 13820 11101 13832 11135
rect 13774 11070 13832 11101
rect 13862 13039 13920 13070
rect 13862 13005 13874 13039
rect 13908 13005 13920 13039
rect 13862 12971 13920 13005
rect 13862 12937 13874 12971
rect 13908 12937 13920 12971
rect 13862 12903 13920 12937
rect 13862 12869 13874 12903
rect 13908 12869 13920 12903
rect 13862 12835 13920 12869
rect 13862 12801 13874 12835
rect 13908 12801 13920 12835
rect 13862 12767 13920 12801
rect 13862 12733 13874 12767
rect 13908 12733 13920 12767
rect 13862 12699 13920 12733
rect 13862 12665 13874 12699
rect 13908 12665 13920 12699
rect 13862 12631 13920 12665
rect 13862 12597 13874 12631
rect 13908 12597 13920 12631
rect 13862 12563 13920 12597
rect 13862 12529 13874 12563
rect 13908 12529 13920 12563
rect 13862 12495 13920 12529
rect 13862 12461 13874 12495
rect 13908 12461 13920 12495
rect 13862 12427 13920 12461
rect 13862 12393 13874 12427
rect 13908 12393 13920 12427
rect 13862 12359 13920 12393
rect 13862 12325 13874 12359
rect 13908 12325 13920 12359
rect 13862 12291 13920 12325
rect 13862 12257 13874 12291
rect 13908 12257 13920 12291
rect 13862 12223 13920 12257
rect 13862 12189 13874 12223
rect 13908 12189 13920 12223
rect 13862 12155 13920 12189
rect 13862 12121 13874 12155
rect 13908 12121 13920 12155
rect 13862 12087 13920 12121
rect 13862 12053 13874 12087
rect 13908 12053 13920 12087
rect 13862 12019 13920 12053
rect 13862 11985 13874 12019
rect 13908 11985 13920 12019
rect 13862 11951 13920 11985
rect 13862 11917 13874 11951
rect 13908 11917 13920 11951
rect 13862 11883 13920 11917
rect 13862 11849 13874 11883
rect 13908 11849 13920 11883
rect 13862 11815 13920 11849
rect 13862 11781 13874 11815
rect 13908 11781 13920 11815
rect 13862 11747 13920 11781
rect 13862 11713 13874 11747
rect 13908 11713 13920 11747
rect 13862 11679 13920 11713
rect 13862 11645 13874 11679
rect 13908 11645 13920 11679
rect 13862 11611 13920 11645
rect 13862 11577 13874 11611
rect 13908 11577 13920 11611
rect 13862 11543 13920 11577
rect 13862 11509 13874 11543
rect 13908 11509 13920 11543
rect 13862 11475 13920 11509
rect 13862 11441 13874 11475
rect 13908 11441 13920 11475
rect 13862 11407 13920 11441
rect 13862 11373 13874 11407
rect 13908 11373 13920 11407
rect 13862 11339 13920 11373
rect 13862 11305 13874 11339
rect 13908 11305 13920 11339
rect 13862 11271 13920 11305
rect 13862 11237 13874 11271
rect 13908 11237 13920 11271
rect 13862 11203 13920 11237
rect 13862 11169 13874 11203
rect 13908 11169 13920 11203
rect 13862 11135 13920 11169
rect 13862 11101 13874 11135
rect 13908 11101 13920 11135
rect 13862 11070 13920 11101
rect 13950 13039 14008 13070
rect 13950 13005 13962 13039
rect 13996 13005 14008 13039
rect 13950 12971 14008 13005
rect 13950 12937 13962 12971
rect 13996 12937 14008 12971
rect 13950 12903 14008 12937
rect 13950 12869 13962 12903
rect 13996 12869 14008 12903
rect 13950 12835 14008 12869
rect 13950 12801 13962 12835
rect 13996 12801 14008 12835
rect 13950 12767 14008 12801
rect 13950 12733 13962 12767
rect 13996 12733 14008 12767
rect 13950 12699 14008 12733
rect 13950 12665 13962 12699
rect 13996 12665 14008 12699
rect 13950 12631 14008 12665
rect 13950 12597 13962 12631
rect 13996 12597 14008 12631
rect 13950 12563 14008 12597
rect 13950 12529 13962 12563
rect 13996 12529 14008 12563
rect 13950 12495 14008 12529
rect 13950 12461 13962 12495
rect 13996 12461 14008 12495
rect 13950 12427 14008 12461
rect 13950 12393 13962 12427
rect 13996 12393 14008 12427
rect 13950 12359 14008 12393
rect 13950 12325 13962 12359
rect 13996 12325 14008 12359
rect 13950 12291 14008 12325
rect 13950 12257 13962 12291
rect 13996 12257 14008 12291
rect 13950 12223 14008 12257
rect 13950 12189 13962 12223
rect 13996 12189 14008 12223
rect 13950 12155 14008 12189
rect 13950 12121 13962 12155
rect 13996 12121 14008 12155
rect 13950 12087 14008 12121
rect 13950 12053 13962 12087
rect 13996 12053 14008 12087
rect 13950 12019 14008 12053
rect 13950 11985 13962 12019
rect 13996 11985 14008 12019
rect 13950 11951 14008 11985
rect 13950 11917 13962 11951
rect 13996 11917 14008 11951
rect 13950 11883 14008 11917
rect 13950 11849 13962 11883
rect 13996 11849 14008 11883
rect 13950 11815 14008 11849
rect 13950 11781 13962 11815
rect 13996 11781 14008 11815
rect 13950 11747 14008 11781
rect 13950 11713 13962 11747
rect 13996 11713 14008 11747
rect 13950 11679 14008 11713
rect 13950 11645 13962 11679
rect 13996 11645 14008 11679
rect 13950 11611 14008 11645
rect 13950 11577 13962 11611
rect 13996 11577 14008 11611
rect 13950 11543 14008 11577
rect 13950 11509 13962 11543
rect 13996 11509 14008 11543
rect 13950 11475 14008 11509
rect 13950 11441 13962 11475
rect 13996 11441 14008 11475
rect 13950 11407 14008 11441
rect 13950 11373 13962 11407
rect 13996 11373 14008 11407
rect 13950 11339 14008 11373
rect 13950 11305 13962 11339
rect 13996 11305 14008 11339
rect 13950 11271 14008 11305
rect 13950 11237 13962 11271
rect 13996 11237 14008 11271
rect 13950 11203 14008 11237
rect 13950 11169 13962 11203
rect 13996 11169 14008 11203
rect 13950 11135 14008 11169
rect 13950 11101 13962 11135
rect 13996 11101 14008 11135
rect 13950 11070 14008 11101
rect 14038 13039 14096 13070
rect 14038 13005 14050 13039
rect 14084 13005 14096 13039
rect 14038 12971 14096 13005
rect 14038 12937 14050 12971
rect 14084 12937 14096 12971
rect 14038 12903 14096 12937
rect 14038 12869 14050 12903
rect 14084 12869 14096 12903
rect 14038 12835 14096 12869
rect 14038 12801 14050 12835
rect 14084 12801 14096 12835
rect 14038 12767 14096 12801
rect 14038 12733 14050 12767
rect 14084 12733 14096 12767
rect 14038 12699 14096 12733
rect 14038 12665 14050 12699
rect 14084 12665 14096 12699
rect 14038 12631 14096 12665
rect 14038 12597 14050 12631
rect 14084 12597 14096 12631
rect 14038 12563 14096 12597
rect 14038 12529 14050 12563
rect 14084 12529 14096 12563
rect 14038 12495 14096 12529
rect 14038 12461 14050 12495
rect 14084 12461 14096 12495
rect 14038 12427 14096 12461
rect 14038 12393 14050 12427
rect 14084 12393 14096 12427
rect 14038 12359 14096 12393
rect 14038 12325 14050 12359
rect 14084 12325 14096 12359
rect 14038 12291 14096 12325
rect 14038 12257 14050 12291
rect 14084 12257 14096 12291
rect 14038 12223 14096 12257
rect 14038 12189 14050 12223
rect 14084 12189 14096 12223
rect 14038 12155 14096 12189
rect 14038 12121 14050 12155
rect 14084 12121 14096 12155
rect 14038 12087 14096 12121
rect 14038 12053 14050 12087
rect 14084 12053 14096 12087
rect 14038 12019 14096 12053
rect 14038 11985 14050 12019
rect 14084 11985 14096 12019
rect 14038 11951 14096 11985
rect 14038 11917 14050 11951
rect 14084 11917 14096 11951
rect 14038 11883 14096 11917
rect 14038 11849 14050 11883
rect 14084 11849 14096 11883
rect 14038 11815 14096 11849
rect 14038 11781 14050 11815
rect 14084 11781 14096 11815
rect 14038 11747 14096 11781
rect 14038 11713 14050 11747
rect 14084 11713 14096 11747
rect 14038 11679 14096 11713
rect 14038 11645 14050 11679
rect 14084 11645 14096 11679
rect 14038 11611 14096 11645
rect 14038 11577 14050 11611
rect 14084 11577 14096 11611
rect 14038 11543 14096 11577
rect 14038 11509 14050 11543
rect 14084 11509 14096 11543
rect 14038 11475 14096 11509
rect 14038 11441 14050 11475
rect 14084 11441 14096 11475
rect 14038 11407 14096 11441
rect 14038 11373 14050 11407
rect 14084 11373 14096 11407
rect 14038 11339 14096 11373
rect 14038 11305 14050 11339
rect 14084 11305 14096 11339
rect 14038 11271 14096 11305
rect 14038 11237 14050 11271
rect 14084 11237 14096 11271
rect 14038 11203 14096 11237
rect 14038 11169 14050 11203
rect 14084 11169 14096 11203
rect 14038 11135 14096 11169
rect 14038 11101 14050 11135
rect 14084 11101 14096 11135
rect 14038 11070 14096 11101
rect 14126 13039 14184 13070
rect 14126 13005 14138 13039
rect 14172 13005 14184 13039
rect 14126 12971 14184 13005
rect 14126 12937 14138 12971
rect 14172 12937 14184 12971
rect 14126 12903 14184 12937
rect 14126 12869 14138 12903
rect 14172 12869 14184 12903
rect 14126 12835 14184 12869
rect 14126 12801 14138 12835
rect 14172 12801 14184 12835
rect 14126 12767 14184 12801
rect 14126 12733 14138 12767
rect 14172 12733 14184 12767
rect 14126 12699 14184 12733
rect 14126 12665 14138 12699
rect 14172 12665 14184 12699
rect 14126 12631 14184 12665
rect 14126 12597 14138 12631
rect 14172 12597 14184 12631
rect 14126 12563 14184 12597
rect 14126 12529 14138 12563
rect 14172 12529 14184 12563
rect 14126 12495 14184 12529
rect 14126 12461 14138 12495
rect 14172 12461 14184 12495
rect 14126 12427 14184 12461
rect 14126 12393 14138 12427
rect 14172 12393 14184 12427
rect 14126 12359 14184 12393
rect 14126 12325 14138 12359
rect 14172 12325 14184 12359
rect 14126 12291 14184 12325
rect 14126 12257 14138 12291
rect 14172 12257 14184 12291
rect 14126 12223 14184 12257
rect 14126 12189 14138 12223
rect 14172 12189 14184 12223
rect 14126 12155 14184 12189
rect 14126 12121 14138 12155
rect 14172 12121 14184 12155
rect 14126 12087 14184 12121
rect 14126 12053 14138 12087
rect 14172 12053 14184 12087
rect 14126 12019 14184 12053
rect 14126 11985 14138 12019
rect 14172 11985 14184 12019
rect 14126 11951 14184 11985
rect 14126 11917 14138 11951
rect 14172 11917 14184 11951
rect 14126 11883 14184 11917
rect 14126 11849 14138 11883
rect 14172 11849 14184 11883
rect 14126 11815 14184 11849
rect 14126 11781 14138 11815
rect 14172 11781 14184 11815
rect 14126 11747 14184 11781
rect 14126 11713 14138 11747
rect 14172 11713 14184 11747
rect 14126 11679 14184 11713
rect 14126 11645 14138 11679
rect 14172 11645 14184 11679
rect 14126 11611 14184 11645
rect 14126 11577 14138 11611
rect 14172 11577 14184 11611
rect 14126 11543 14184 11577
rect 14126 11509 14138 11543
rect 14172 11509 14184 11543
rect 14126 11475 14184 11509
rect 14126 11441 14138 11475
rect 14172 11441 14184 11475
rect 14126 11407 14184 11441
rect 14126 11373 14138 11407
rect 14172 11373 14184 11407
rect 14126 11339 14184 11373
rect 14126 11305 14138 11339
rect 14172 11305 14184 11339
rect 14126 11271 14184 11305
rect 14126 11237 14138 11271
rect 14172 11237 14184 11271
rect 14126 11203 14184 11237
rect 14126 11169 14138 11203
rect 14172 11169 14184 11203
rect 14126 11135 14184 11169
rect 14126 11101 14138 11135
rect 14172 11101 14184 11135
rect 14126 11070 14184 11101
rect 14214 13039 14272 13070
rect 14214 13005 14226 13039
rect 14260 13005 14272 13039
rect 14214 12971 14272 13005
rect 14214 12937 14226 12971
rect 14260 12937 14272 12971
rect 14214 12903 14272 12937
rect 14214 12869 14226 12903
rect 14260 12869 14272 12903
rect 14214 12835 14272 12869
rect 14214 12801 14226 12835
rect 14260 12801 14272 12835
rect 14214 12767 14272 12801
rect 14214 12733 14226 12767
rect 14260 12733 14272 12767
rect 14214 12699 14272 12733
rect 14214 12665 14226 12699
rect 14260 12665 14272 12699
rect 14214 12631 14272 12665
rect 14214 12597 14226 12631
rect 14260 12597 14272 12631
rect 14214 12563 14272 12597
rect 14214 12529 14226 12563
rect 14260 12529 14272 12563
rect 14214 12495 14272 12529
rect 14214 12461 14226 12495
rect 14260 12461 14272 12495
rect 14214 12427 14272 12461
rect 14214 12393 14226 12427
rect 14260 12393 14272 12427
rect 14214 12359 14272 12393
rect 14214 12325 14226 12359
rect 14260 12325 14272 12359
rect 14214 12291 14272 12325
rect 14214 12257 14226 12291
rect 14260 12257 14272 12291
rect 14214 12223 14272 12257
rect 14214 12189 14226 12223
rect 14260 12189 14272 12223
rect 14214 12155 14272 12189
rect 14214 12121 14226 12155
rect 14260 12121 14272 12155
rect 14214 12087 14272 12121
rect 14214 12053 14226 12087
rect 14260 12053 14272 12087
rect 14214 12019 14272 12053
rect 14214 11985 14226 12019
rect 14260 11985 14272 12019
rect 14214 11951 14272 11985
rect 14214 11917 14226 11951
rect 14260 11917 14272 11951
rect 14214 11883 14272 11917
rect 14214 11849 14226 11883
rect 14260 11849 14272 11883
rect 14214 11815 14272 11849
rect 14214 11781 14226 11815
rect 14260 11781 14272 11815
rect 14214 11747 14272 11781
rect 14214 11713 14226 11747
rect 14260 11713 14272 11747
rect 14214 11679 14272 11713
rect 14214 11645 14226 11679
rect 14260 11645 14272 11679
rect 14214 11611 14272 11645
rect 14214 11577 14226 11611
rect 14260 11577 14272 11611
rect 14214 11543 14272 11577
rect 14214 11509 14226 11543
rect 14260 11509 14272 11543
rect 14214 11475 14272 11509
rect 14214 11441 14226 11475
rect 14260 11441 14272 11475
rect 14214 11407 14272 11441
rect 14214 11373 14226 11407
rect 14260 11373 14272 11407
rect 14214 11339 14272 11373
rect 14214 11305 14226 11339
rect 14260 11305 14272 11339
rect 14214 11271 14272 11305
rect 14214 11237 14226 11271
rect 14260 11237 14272 11271
rect 14214 11203 14272 11237
rect 14214 11169 14226 11203
rect 14260 11169 14272 11203
rect 14214 11135 14272 11169
rect 14214 11101 14226 11135
rect 14260 11101 14272 11135
rect 14214 11070 14272 11101
rect 14302 13039 14360 13070
rect 14302 13005 14314 13039
rect 14348 13005 14360 13039
rect 14302 12971 14360 13005
rect 14302 12937 14314 12971
rect 14348 12937 14360 12971
rect 14302 12903 14360 12937
rect 14302 12869 14314 12903
rect 14348 12869 14360 12903
rect 14302 12835 14360 12869
rect 14302 12801 14314 12835
rect 14348 12801 14360 12835
rect 14302 12767 14360 12801
rect 14302 12733 14314 12767
rect 14348 12733 14360 12767
rect 14302 12699 14360 12733
rect 14302 12665 14314 12699
rect 14348 12665 14360 12699
rect 14302 12631 14360 12665
rect 14302 12597 14314 12631
rect 14348 12597 14360 12631
rect 14302 12563 14360 12597
rect 14302 12529 14314 12563
rect 14348 12529 14360 12563
rect 14302 12495 14360 12529
rect 14302 12461 14314 12495
rect 14348 12461 14360 12495
rect 14302 12427 14360 12461
rect 14302 12393 14314 12427
rect 14348 12393 14360 12427
rect 14302 12359 14360 12393
rect 14302 12325 14314 12359
rect 14348 12325 14360 12359
rect 14302 12291 14360 12325
rect 14302 12257 14314 12291
rect 14348 12257 14360 12291
rect 14302 12223 14360 12257
rect 14302 12189 14314 12223
rect 14348 12189 14360 12223
rect 14302 12155 14360 12189
rect 14302 12121 14314 12155
rect 14348 12121 14360 12155
rect 14302 12087 14360 12121
rect 14302 12053 14314 12087
rect 14348 12053 14360 12087
rect 14302 12019 14360 12053
rect 14302 11985 14314 12019
rect 14348 11985 14360 12019
rect 14302 11951 14360 11985
rect 14302 11917 14314 11951
rect 14348 11917 14360 11951
rect 14302 11883 14360 11917
rect 14302 11849 14314 11883
rect 14348 11849 14360 11883
rect 14302 11815 14360 11849
rect 14302 11781 14314 11815
rect 14348 11781 14360 11815
rect 14302 11747 14360 11781
rect 14302 11713 14314 11747
rect 14348 11713 14360 11747
rect 14302 11679 14360 11713
rect 14302 11645 14314 11679
rect 14348 11645 14360 11679
rect 14302 11611 14360 11645
rect 14302 11577 14314 11611
rect 14348 11577 14360 11611
rect 14302 11543 14360 11577
rect 14302 11509 14314 11543
rect 14348 11509 14360 11543
rect 14302 11475 14360 11509
rect 14302 11441 14314 11475
rect 14348 11441 14360 11475
rect 14302 11407 14360 11441
rect 14302 11373 14314 11407
rect 14348 11373 14360 11407
rect 14302 11339 14360 11373
rect 14302 11305 14314 11339
rect 14348 11305 14360 11339
rect 14302 11271 14360 11305
rect 14302 11237 14314 11271
rect 14348 11237 14360 11271
rect 14302 11203 14360 11237
rect 14302 11169 14314 11203
rect 14348 11169 14360 11203
rect 14302 11135 14360 11169
rect 14302 11101 14314 11135
rect 14348 11101 14360 11135
rect 14302 11070 14360 11101
rect 14390 13039 14448 13070
rect 14390 13005 14402 13039
rect 14436 13005 14448 13039
rect 14390 12971 14448 13005
rect 14390 12937 14402 12971
rect 14436 12937 14448 12971
rect 14390 12903 14448 12937
rect 14390 12869 14402 12903
rect 14436 12869 14448 12903
rect 14390 12835 14448 12869
rect 14390 12801 14402 12835
rect 14436 12801 14448 12835
rect 14390 12767 14448 12801
rect 14390 12733 14402 12767
rect 14436 12733 14448 12767
rect 14390 12699 14448 12733
rect 14390 12665 14402 12699
rect 14436 12665 14448 12699
rect 14390 12631 14448 12665
rect 14390 12597 14402 12631
rect 14436 12597 14448 12631
rect 14390 12563 14448 12597
rect 14390 12529 14402 12563
rect 14436 12529 14448 12563
rect 14390 12495 14448 12529
rect 14390 12461 14402 12495
rect 14436 12461 14448 12495
rect 14390 12427 14448 12461
rect 14390 12393 14402 12427
rect 14436 12393 14448 12427
rect 14390 12359 14448 12393
rect 14390 12325 14402 12359
rect 14436 12325 14448 12359
rect 14390 12291 14448 12325
rect 14390 12257 14402 12291
rect 14436 12257 14448 12291
rect 14390 12223 14448 12257
rect 14390 12189 14402 12223
rect 14436 12189 14448 12223
rect 14390 12155 14448 12189
rect 14390 12121 14402 12155
rect 14436 12121 14448 12155
rect 14390 12087 14448 12121
rect 14390 12053 14402 12087
rect 14436 12053 14448 12087
rect 14390 12019 14448 12053
rect 14390 11985 14402 12019
rect 14436 11985 14448 12019
rect 14390 11951 14448 11985
rect 14390 11917 14402 11951
rect 14436 11917 14448 11951
rect 14390 11883 14448 11917
rect 14390 11849 14402 11883
rect 14436 11849 14448 11883
rect 14390 11815 14448 11849
rect 14390 11781 14402 11815
rect 14436 11781 14448 11815
rect 14390 11747 14448 11781
rect 14390 11713 14402 11747
rect 14436 11713 14448 11747
rect 14390 11679 14448 11713
rect 14390 11645 14402 11679
rect 14436 11645 14448 11679
rect 14390 11611 14448 11645
rect 14390 11577 14402 11611
rect 14436 11577 14448 11611
rect 14390 11543 14448 11577
rect 14390 11509 14402 11543
rect 14436 11509 14448 11543
rect 14390 11475 14448 11509
rect 14390 11441 14402 11475
rect 14436 11441 14448 11475
rect 14390 11407 14448 11441
rect 14390 11373 14402 11407
rect 14436 11373 14448 11407
rect 14390 11339 14448 11373
rect 14390 11305 14402 11339
rect 14436 11305 14448 11339
rect 14390 11271 14448 11305
rect 14390 11237 14402 11271
rect 14436 11237 14448 11271
rect 14390 11203 14448 11237
rect 14390 11169 14402 11203
rect 14436 11169 14448 11203
rect 14390 11135 14448 11169
rect 14390 11101 14402 11135
rect 14436 11101 14448 11135
rect 14390 11070 14448 11101
rect 14478 13039 14536 13070
rect 14478 13005 14490 13039
rect 14524 13005 14536 13039
rect 14478 12971 14536 13005
rect 14478 12937 14490 12971
rect 14524 12937 14536 12971
rect 14478 12903 14536 12937
rect 14478 12869 14490 12903
rect 14524 12869 14536 12903
rect 14478 12835 14536 12869
rect 14478 12801 14490 12835
rect 14524 12801 14536 12835
rect 14478 12767 14536 12801
rect 14478 12733 14490 12767
rect 14524 12733 14536 12767
rect 14478 12699 14536 12733
rect 14478 12665 14490 12699
rect 14524 12665 14536 12699
rect 14478 12631 14536 12665
rect 14478 12597 14490 12631
rect 14524 12597 14536 12631
rect 14478 12563 14536 12597
rect 14478 12529 14490 12563
rect 14524 12529 14536 12563
rect 14478 12495 14536 12529
rect 14478 12461 14490 12495
rect 14524 12461 14536 12495
rect 14478 12427 14536 12461
rect 14478 12393 14490 12427
rect 14524 12393 14536 12427
rect 14478 12359 14536 12393
rect 14478 12325 14490 12359
rect 14524 12325 14536 12359
rect 14478 12291 14536 12325
rect 14478 12257 14490 12291
rect 14524 12257 14536 12291
rect 14478 12223 14536 12257
rect 14478 12189 14490 12223
rect 14524 12189 14536 12223
rect 14478 12155 14536 12189
rect 14478 12121 14490 12155
rect 14524 12121 14536 12155
rect 14478 12087 14536 12121
rect 14478 12053 14490 12087
rect 14524 12053 14536 12087
rect 14478 12019 14536 12053
rect 14478 11985 14490 12019
rect 14524 11985 14536 12019
rect 14478 11951 14536 11985
rect 14478 11917 14490 11951
rect 14524 11917 14536 11951
rect 14478 11883 14536 11917
rect 14478 11849 14490 11883
rect 14524 11849 14536 11883
rect 14478 11815 14536 11849
rect 14478 11781 14490 11815
rect 14524 11781 14536 11815
rect 14478 11747 14536 11781
rect 14478 11713 14490 11747
rect 14524 11713 14536 11747
rect 14478 11679 14536 11713
rect 14478 11645 14490 11679
rect 14524 11645 14536 11679
rect 14478 11611 14536 11645
rect 14478 11577 14490 11611
rect 14524 11577 14536 11611
rect 14478 11543 14536 11577
rect 14478 11509 14490 11543
rect 14524 11509 14536 11543
rect 14478 11475 14536 11509
rect 14478 11441 14490 11475
rect 14524 11441 14536 11475
rect 14478 11407 14536 11441
rect 14478 11373 14490 11407
rect 14524 11373 14536 11407
rect 14478 11339 14536 11373
rect 14478 11305 14490 11339
rect 14524 11305 14536 11339
rect 14478 11271 14536 11305
rect 14478 11237 14490 11271
rect 14524 11237 14536 11271
rect 14478 11203 14536 11237
rect 14478 11169 14490 11203
rect 14524 11169 14536 11203
rect 14478 11135 14536 11169
rect 14478 11101 14490 11135
rect 14524 11101 14536 11135
rect 14478 11070 14536 11101
rect 14566 13039 14624 13070
rect 14566 13005 14578 13039
rect 14612 13005 14624 13039
rect 14566 12971 14624 13005
rect 14566 12937 14578 12971
rect 14612 12937 14624 12971
rect 14566 12903 14624 12937
rect 14566 12869 14578 12903
rect 14612 12869 14624 12903
rect 14566 12835 14624 12869
rect 14566 12801 14578 12835
rect 14612 12801 14624 12835
rect 14566 12767 14624 12801
rect 14566 12733 14578 12767
rect 14612 12733 14624 12767
rect 14566 12699 14624 12733
rect 14566 12665 14578 12699
rect 14612 12665 14624 12699
rect 14566 12631 14624 12665
rect 14566 12597 14578 12631
rect 14612 12597 14624 12631
rect 14566 12563 14624 12597
rect 14566 12529 14578 12563
rect 14612 12529 14624 12563
rect 14566 12495 14624 12529
rect 14566 12461 14578 12495
rect 14612 12461 14624 12495
rect 14566 12427 14624 12461
rect 14566 12393 14578 12427
rect 14612 12393 14624 12427
rect 14566 12359 14624 12393
rect 14566 12325 14578 12359
rect 14612 12325 14624 12359
rect 14566 12291 14624 12325
rect 14566 12257 14578 12291
rect 14612 12257 14624 12291
rect 14566 12223 14624 12257
rect 14566 12189 14578 12223
rect 14612 12189 14624 12223
rect 14566 12155 14624 12189
rect 14566 12121 14578 12155
rect 14612 12121 14624 12155
rect 14566 12087 14624 12121
rect 14566 12053 14578 12087
rect 14612 12053 14624 12087
rect 14566 12019 14624 12053
rect 14566 11985 14578 12019
rect 14612 11985 14624 12019
rect 14566 11951 14624 11985
rect 14566 11917 14578 11951
rect 14612 11917 14624 11951
rect 14566 11883 14624 11917
rect 14566 11849 14578 11883
rect 14612 11849 14624 11883
rect 14566 11815 14624 11849
rect 14566 11781 14578 11815
rect 14612 11781 14624 11815
rect 14566 11747 14624 11781
rect 14566 11713 14578 11747
rect 14612 11713 14624 11747
rect 14566 11679 14624 11713
rect 14566 11645 14578 11679
rect 14612 11645 14624 11679
rect 14566 11611 14624 11645
rect 14566 11577 14578 11611
rect 14612 11577 14624 11611
rect 14566 11543 14624 11577
rect 14566 11509 14578 11543
rect 14612 11509 14624 11543
rect 14566 11475 14624 11509
rect 14566 11441 14578 11475
rect 14612 11441 14624 11475
rect 14566 11407 14624 11441
rect 14566 11373 14578 11407
rect 14612 11373 14624 11407
rect 14566 11339 14624 11373
rect 14566 11305 14578 11339
rect 14612 11305 14624 11339
rect 14566 11271 14624 11305
rect 14566 11237 14578 11271
rect 14612 11237 14624 11271
rect 14566 11203 14624 11237
rect 14566 11169 14578 11203
rect 14612 11169 14624 11203
rect 14566 11135 14624 11169
rect 14566 11101 14578 11135
rect 14612 11101 14624 11135
rect 14566 11070 14624 11101
rect 14654 13039 14712 13070
rect 14654 13005 14666 13039
rect 14700 13005 14712 13039
rect 14654 12971 14712 13005
rect 14654 12937 14666 12971
rect 14700 12937 14712 12971
rect 14654 12903 14712 12937
rect 14654 12869 14666 12903
rect 14700 12869 14712 12903
rect 14654 12835 14712 12869
rect 14654 12801 14666 12835
rect 14700 12801 14712 12835
rect 14654 12767 14712 12801
rect 14654 12733 14666 12767
rect 14700 12733 14712 12767
rect 14654 12699 14712 12733
rect 14654 12665 14666 12699
rect 14700 12665 14712 12699
rect 14654 12631 14712 12665
rect 14654 12597 14666 12631
rect 14700 12597 14712 12631
rect 14654 12563 14712 12597
rect 14654 12529 14666 12563
rect 14700 12529 14712 12563
rect 14654 12495 14712 12529
rect 14654 12461 14666 12495
rect 14700 12461 14712 12495
rect 14654 12427 14712 12461
rect 14654 12393 14666 12427
rect 14700 12393 14712 12427
rect 14654 12359 14712 12393
rect 14654 12325 14666 12359
rect 14700 12325 14712 12359
rect 14654 12291 14712 12325
rect 14654 12257 14666 12291
rect 14700 12257 14712 12291
rect 14654 12223 14712 12257
rect 14654 12189 14666 12223
rect 14700 12189 14712 12223
rect 14654 12155 14712 12189
rect 14654 12121 14666 12155
rect 14700 12121 14712 12155
rect 14654 12087 14712 12121
rect 14654 12053 14666 12087
rect 14700 12053 14712 12087
rect 14654 12019 14712 12053
rect 14654 11985 14666 12019
rect 14700 11985 14712 12019
rect 14654 11951 14712 11985
rect 14654 11917 14666 11951
rect 14700 11917 14712 11951
rect 14654 11883 14712 11917
rect 14654 11849 14666 11883
rect 14700 11849 14712 11883
rect 14654 11815 14712 11849
rect 14654 11781 14666 11815
rect 14700 11781 14712 11815
rect 14654 11747 14712 11781
rect 14654 11713 14666 11747
rect 14700 11713 14712 11747
rect 14654 11679 14712 11713
rect 14654 11645 14666 11679
rect 14700 11645 14712 11679
rect 14654 11611 14712 11645
rect 14654 11577 14666 11611
rect 14700 11577 14712 11611
rect 14654 11543 14712 11577
rect 14654 11509 14666 11543
rect 14700 11509 14712 11543
rect 14654 11475 14712 11509
rect 14654 11441 14666 11475
rect 14700 11441 14712 11475
rect 14654 11407 14712 11441
rect 14654 11373 14666 11407
rect 14700 11373 14712 11407
rect 14654 11339 14712 11373
rect 14654 11305 14666 11339
rect 14700 11305 14712 11339
rect 14654 11271 14712 11305
rect 14654 11237 14666 11271
rect 14700 11237 14712 11271
rect 14654 11203 14712 11237
rect 14654 11169 14666 11203
rect 14700 11169 14712 11203
rect 14654 11135 14712 11169
rect 14654 11101 14666 11135
rect 14700 11101 14712 11135
rect 14654 11070 14712 11101
rect 14742 13039 14800 13070
rect 14742 13005 14754 13039
rect 14788 13005 14800 13039
rect 14742 12971 14800 13005
rect 14742 12937 14754 12971
rect 14788 12937 14800 12971
rect 14742 12903 14800 12937
rect 14742 12869 14754 12903
rect 14788 12869 14800 12903
rect 14742 12835 14800 12869
rect 14742 12801 14754 12835
rect 14788 12801 14800 12835
rect 14742 12767 14800 12801
rect 14742 12733 14754 12767
rect 14788 12733 14800 12767
rect 14742 12699 14800 12733
rect 14742 12665 14754 12699
rect 14788 12665 14800 12699
rect 14742 12631 14800 12665
rect 14742 12597 14754 12631
rect 14788 12597 14800 12631
rect 14742 12563 14800 12597
rect 14742 12529 14754 12563
rect 14788 12529 14800 12563
rect 14742 12495 14800 12529
rect 14742 12461 14754 12495
rect 14788 12461 14800 12495
rect 14742 12427 14800 12461
rect 14742 12393 14754 12427
rect 14788 12393 14800 12427
rect 14742 12359 14800 12393
rect 14742 12325 14754 12359
rect 14788 12325 14800 12359
rect 14742 12291 14800 12325
rect 14742 12257 14754 12291
rect 14788 12257 14800 12291
rect 14742 12223 14800 12257
rect 14742 12189 14754 12223
rect 14788 12189 14800 12223
rect 14742 12155 14800 12189
rect 14742 12121 14754 12155
rect 14788 12121 14800 12155
rect 14742 12087 14800 12121
rect 14742 12053 14754 12087
rect 14788 12053 14800 12087
rect 14742 12019 14800 12053
rect 14742 11985 14754 12019
rect 14788 11985 14800 12019
rect 14742 11951 14800 11985
rect 14742 11917 14754 11951
rect 14788 11917 14800 11951
rect 14742 11883 14800 11917
rect 14742 11849 14754 11883
rect 14788 11849 14800 11883
rect 14742 11815 14800 11849
rect 14742 11781 14754 11815
rect 14788 11781 14800 11815
rect 14742 11747 14800 11781
rect 14742 11713 14754 11747
rect 14788 11713 14800 11747
rect 14742 11679 14800 11713
rect 14742 11645 14754 11679
rect 14788 11645 14800 11679
rect 14742 11611 14800 11645
rect 14742 11577 14754 11611
rect 14788 11577 14800 11611
rect 14742 11543 14800 11577
rect 14742 11509 14754 11543
rect 14788 11509 14800 11543
rect 14742 11475 14800 11509
rect 14742 11441 14754 11475
rect 14788 11441 14800 11475
rect 14742 11407 14800 11441
rect 14742 11373 14754 11407
rect 14788 11373 14800 11407
rect 14742 11339 14800 11373
rect 14742 11305 14754 11339
rect 14788 11305 14800 11339
rect 14742 11271 14800 11305
rect 14742 11237 14754 11271
rect 14788 11237 14800 11271
rect 14742 11203 14800 11237
rect 14742 11169 14754 11203
rect 14788 11169 14800 11203
rect 14742 11135 14800 11169
rect 14742 11101 14754 11135
rect 14788 11101 14800 11135
rect 14742 11070 14800 11101
rect 14830 13039 14888 13070
rect 14830 13005 14842 13039
rect 14876 13005 14888 13039
rect 14830 12971 14888 13005
rect 14830 12937 14842 12971
rect 14876 12937 14888 12971
rect 14830 12903 14888 12937
rect 14830 12869 14842 12903
rect 14876 12869 14888 12903
rect 14830 12835 14888 12869
rect 14830 12801 14842 12835
rect 14876 12801 14888 12835
rect 14830 12767 14888 12801
rect 14830 12733 14842 12767
rect 14876 12733 14888 12767
rect 14830 12699 14888 12733
rect 14830 12665 14842 12699
rect 14876 12665 14888 12699
rect 14830 12631 14888 12665
rect 14830 12597 14842 12631
rect 14876 12597 14888 12631
rect 14830 12563 14888 12597
rect 14830 12529 14842 12563
rect 14876 12529 14888 12563
rect 14830 12495 14888 12529
rect 14830 12461 14842 12495
rect 14876 12461 14888 12495
rect 14830 12427 14888 12461
rect 14830 12393 14842 12427
rect 14876 12393 14888 12427
rect 14830 12359 14888 12393
rect 14830 12325 14842 12359
rect 14876 12325 14888 12359
rect 14830 12291 14888 12325
rect 14830 12257 14842 12291
rect 14876 12257 14888 12291
rect 14830 12223 14888 12257
rect 14830 12189 14842 12223
rect 14876 12189 14888 12223
rect 14830 12155 14888 12189
rect 14830 12121 14842 12155
rect 14876 12121 14888 12155
rect 14830 12087 14888 12121
rect 14830 12053 14842 12087
rect 14876 12053 14888 12087
rect 14830 12019 14888 12053
rect 14830 11985 14842 12019
rect 14876 11985 14888 12019
rect 14830 11951 14888 11985
rect 14830 11917 14842 11951
rect 14876 11917 14888 11951
rect 14830 11883 14888 11917
rect 14830 11849 14842 11883
rect 14876 11849 14888 11883
rect 14830 11815 14888 11849
rect 14830 11781 14842 11815
rect 14876 11781 14888 11815
rect 14830 11747 14888 11781
rect 14830 11713 14842 11747
rect 14876 11713 14888 11747
rect 14830 11679 14888 11713
rect 14830 11645 14842 11679
rect 14876 11645 14888 11679
rect 14830 11611 14888 11645
rect 14830 11577 14842 11611
rect 14876 11577 14888 11611
rect 14830 11543 14888 11577
rect 14830 11509 14842 11543
rect 14876 11509 14888 11543
rect 14830 11475 14888 11509
rect 14830 11441 14842 11475
rect 14876 11441 14888 11475
rect 14830 11407 14888 11441
rect 14830 11373 14842 11407
rect 14876 11373 14888 11407
rect 14830 11339 14888 11373
rect 14830 11305 14842 11339
rect 14876 11305 14888 11339
rect 14830 11271 14888 11305
rect 14830 11237 14842 11271
rect 14876 11237 14888 11271
rect 14830 11203 14888 11237
rect 14830 11169 14842 11203
rect 14876 11169 14888 11203
rect 14830 11135 14888 11169
rect 14830 11101 14842 11135
rect 14876 11101 14888 11135
rect 14830 11070 14888 11101
rect 14918 13039 14976 13070
rect 14918 13005 14930 13039
rect 14964 13005 14976 13039
rect 14918 12971 14976 13005
rect 14918 12937 14930 12971
rect 14964 12937 14976 12971
rect 14918 12903 14976 12937
rect 14918 12869 14930 12903
rect 14964 12869 14976 12903
rect 14918 12835 14976 12869
rect 14918 12801 14930 12835
rect 14964 12801 14976 12835
rect 14918 12767 14976 12801
rect 14918 12733 14930 12767
rect 14964 12733 14976 12767
rect 14918 12699 14976 12733
rect 14918 12665 14930 12699
rect 14964 12665 14976 12699
rect 14918 12631 14976 12665
rect 14918 12597 14930 12631
rect 14964 12597 14976 12631
rect 14918 12563 14976 12597
rect 14918 12529 14930 12563
rect 14964 12529 14976 12563
rect 14918 12495 14976 12529
rect 14918 12461 14930 12495
rect 14964 12461 14976 12495
rect 14918 12427 14976 12461
rect 14918 12393 14930 12427
rect 14964 12393 14976 12427
rect 14918 12359 14976 12393
rect 14918 12325 14930 12359
rect 14964 12325 14976 12359
rect 14918 12291 14976 12325
rect 14918 12257 14930 12291
rect 14964 12257 14976 12291
rect 14918 12223 14976 12257
rect 14918 12189 14930 12223
rect 14964 12189 14976 12223
rect 14918 12155 14976 12189
rect 14918 12121 14930 12155
rect 14964 12121 14976 12155
rect 14918 12087 14976 12121
rect 14918 12053 14930 12087
rect 14964 12053 14976 12087
rect 14918 12019 14976 12053
rect 14918 11985 14930 12019
rect 14964 11985 14976 12019
rect 14918 11951 14976 11985
rect 14918 11917 14930 11951
rect 14964 11917 14976 11951
rect 14918 11883 14976 11917
rect 14918 11849 14930 11883
rect 14964 11849 14976 11883
rect 14918 11815 14976 11849
rect 14918 11781 14930 11815
rect 14964 11781 14976 11815
rect 14918 11747 14976 11781
rect 14918 11713 14930 11747
rect 14964 11713 14976 11747
rect 14918 11679 14976 11713
rect 14918 11645 14930 11679
rect 14964 11645 14976 11679
rect 14918 11611 14976 11645
rect 14918 11577 14930 11611
rect 14964 11577 14976 11611
rect 14918 11543 14976 11577
rect 14918 11509 14930 11543
rect 14964 11509 14976 11543
rect 14918 11475 14976 11509
rect 14918 11441 14930 11475
rect 14964 11441 14976 11475
rect 14918 11407 14976 11441
rect 14918 11373 14930 11407
rect 14964 11373 14976 11407
rect 14918 11339 14976 11373
rect 14918 11305 14930 11339
rect 14964 11305 14976 11339
rect 14918 11271 14976 11305
rect 14918 11237 14930 11271
rect 14964 11237 14976 11271
rect 14918 11203 14976 11237
rect 14918 11169 14930 11203
rect 14964 11169 14976 11203
rect 14918 11135 14976 11169
rect 14918 11101 14930 11135
rect 14964 11101 14976 11135
rect 14918 11070 14976 11101
rect 15006 13039 15064 13070
rect 15006 13005 15018 13039
rect 15052 13005 15064 13039
rect 15006 12971 15064 13005
rect 15006 12937 15018 12971
rect 15052 12937 15064 12971
rect 15006 12903 15064 12937
rect 15006 12869 15018 12903
rect 15052 12869 15064 12903
rect 15006 12835 15064 12869
rect 15006 12801 15018 12835
rect 15052 12801 15064 12835
rect 15006 12767 15064 12801
rect 15006 12733 15018 12767
rect 15052 12733 15064 12767
rect 15006 12699 15064 12733
rect 15006 12665 15018 12699
rect 15052 12665 15064 12699
rect 15006 12631 15064 12665
rect 15006 12597 15018 12631
rect 15052 12597 15064 12631
rect 15006 12563 15064 12597
rect 15006 12529 15018 12563
rect 15052 12529 15064 12563
rect 15006 12495 15064 12529
rect 15006 12461 15018 12495
rect 15052 12461 15064 12495
rect 15006 12427 15064 12461
rect 15006 12393 15018 12427
rect 15052 12393 15064 12427
rect 15006 12359 15064 12393
rect 15006 12325 15018 12359
rect 15052 12325 15064 12359
rect 15006 12291 15064 12325
rect 15006 12257 15018 12291
rect 15052 12257 15064 12291
rect 15006 12223 15064 12257
rect 15006 12189 15018 12223
rect 15052 12189 15064 12223
rect 15006 12155 15064 12189
rect 15006 12121 15018 12155
rect 15052 12121 15064 12155
rect 15006 12087 15064 12121
rect 15006 12053 15018 12087
rect 15052 12053 15064 12087
rect 15006 12019 15064 12053
rect 15006 11985 15018 12019
rect 15052 11985 15064 12019
rect 15006 11951 15064 11985
rect 15006 11917 15018 11951
rect 15052 11917 15064 11951
rect 15006 11883 15064 11917
rect 15006 11849 15018 11883
rect 15052 11849 15064 11883
rect 15006 11815 15064 11849
rect 15006 11781 15018 11815
rect 15052 11781 15064 11815
rect 15006 11747 15064 11781
rect 15006 11713 15018 11747
rect 15052 11713 15064 11747
rect 15006 11679 15064 11713
rect 15006 11645 15018 11679
rect 15052 11645 15064 11679
rect 15006 11611 15064 11645
rect 15006 11577 15018 11611
rect 15052 11577 15064 11611
rect 15006 11543 15064 11577
rect 15006 11509 15018 11543
rect 15052 11509 15064 11543
rect 15006 11475 15064 11509
rect 15006 11441 15018 11475
rect 15052 11441 15064 11475
rect 15006 11407 15064 11441
rect 15006 11373 15018 11407
rect 15052 11373 15064 11407
rect 15006 11339 15064 11373
rect 15006 11305 15018 11339
rect 15052 11305 15064 11339
rect 15006 11271 15064 11305
rect 15006 11237 15018 11271
rect 15052 11237 15064 11271
rect 15006 11203 15064 11237
rect 15006 11169 15018 11203
rect 15052 11169 15064 11203
rect 15006 11135 15064 11169
rect 15006 11101 15018 11135
rect 15052 11101 15064 11135
rect 15006 11070 15064 11101
rect 15094 13039 15152 13070
rect 15094 13005 15106 13039
rect 15140 13005 15152 13039
rect 15094 12971 15152 13005
rect 15094 12937 15106 12971
rect 15140 12937 15152 12971
rect 15094 12903 15152 12937
rect 15094 12869 15106 12903
rect 15140 12869 15152 12903
rect 15094 12835 15152 12869
rect 15094 12801 15106 12835
rect 15140 12801 15152 12835
rect 15094 12767 15152 12801
rect 15094 12733 15106 12767
rect 15140 12733 15152 12767
rect 15094 12699 15152 12733
rect 15094 12665 15106 12699
rect 15140 12665 15152 12699
rect 15094 12631 15152 12665
rect 15094 12597 15106 12631
rect 15140 12597 15152 12631
rect 15094 12563 15152 12597
rect 15094 12529 15106 12563
rect 15140 12529 15152 12563
rect 15094 12495 15152 12529
rect 15094 12461 15106 12495
rect 15140 12461 15152 12495
rect 15094 12427 15152 12461
rect 15094 12393 15106 12427
rect 15140 12393 15152 12427
rect 15094 12359 15152 12393
rect 15094 12325 15106 12359
rect 15140 12325 15152 12359
rect 15094 12291 15152 12325
rect 15094 12257 15106 12291
rect 15140 12257 15152 12291
rect 15094 12223 15152 12257
rect 15094 12189 15106 12223
rect 15140 12189 15152 12223
rect 15094 12155 15152 12189
rect 15094 12121 15106 12155
rect 15140 12121 15152 12155
rect 15094 12087 15152 12121
rect 15094 12053 15106 12087
rect 15140 12053 15152 12087
rect 15094 12019 15152 12053
rect 15094 11985 15106 12019
rect 15140 11985 15152 12019
rect 15094 11951 15152 11985
rect 15094 11917 15106 11951
rect 15140 11917 15152 11951
rect 15094 11883 15152 11917
rect 15094 11849 15106 11883
rect 15140 11849 15152 11883
rect 15094 11815 15152 11849
rect 15094 11781 15106 11815
rect 15140 11781 15152 11815
rect 15094 11747 15152 11781
rect 15094 11713 15106 11747
rect 15140 11713 15152 11747
rect 15094 11679 15152 11713
rect 15094 11645 15106 11679
rect 15140 11645 15152 11679
rect 15094 11611 15152 11645
rect 15094 11577 15106 11611
rect 15140 11577 15152 11611
rect 15094 11543 15152 11577
rect 15094 11509 15106 11543
rect 15140 11509 15152 11543
rect 15094 11475 15152 11509
rect 15094 11441 15106 11475
rect 15140 11441 15152 11475
rect 15094 11407 15152 11441
rect 15094 11373 15106 11407
rect 15140 11373 15152 11407
rect 15094 11339 15152 11373
rect 15094 11305 15106 11339
rect 15140 11305 15152 11339
rect 15094 11271 15152 11305
rect 15094 11237 15106 11271
rect 15140 11237 15152 11271
rect 15094 11203 15152 11237
rect 15094 11169 15106 11203
rect 15140 11169 15152 11203
rect 15094 11135 15152 11169
rect 15094 11101 15106 11135
rect 15140 11101 15152 11135
rect 15094 11070 15152 11101
rect 15182 13039 15240 13070
rect 15182 13005 15194 13039
rect 15228 13005 15240 13039
rect 15182 12971 15240 13005
rect 15182 12937 15194 12971
rect 15228 12937 15240 12971
rect 15182 12903 15240 12937
rect 15182 12869 15194 12903
rect 15228 12869 15240 12903
rect 15182 12835 15240 12869
rect 15182 12801 15194 12835
rect 15228 12801 15240 12835
rect 15182 12767 15240 12801
rect 15182 12733 15194 12767
rect 15228 12733 15240 12767
rect 15182 12699 15240 12733
rect 15182 12665 15194 12699
rect 15228 12665 15240 12699
rect 15182 12631 15240 12665
rect 15182 12597 15194 12631
rect 15228 12597 15240 12631
rect 15182 12563 15240 12597
rect 15182 12529 15194 12563
rect 15228 12529 15240 12563
rect 15182 12495 15240 12529
rect 15182 12461 15194 12495
rect 15228 12461 15240 12495
rect 15182 12427 15240 12461
rect 15182 12393 15194 12427
rect 15228 12393 15240 12427
rect 15182 12359 15240 12393
rect 15182 12325 15194 12359
rect 15228 12325 15240 12359
rect 15182 12291 15240 12325
rect 15182 12257 15194 12291
rect 15228 12257 15240 12291
rect 15182 12223 15240 12257
rect 15182 12189 15194 12223
rect 15228 12189 15240 12223
rect 15182 12155 15240 12189
rect 15182 12121 15194 12155
rect 15228 12121 15240 12155
rect 15182 12087 15240 12121
rect 15182 12053 15194 12087
rect 15228 12053 15240 12087
rect 15182 12019 15240 12053
rect 15182 11985 15194 12019
rect 15228 11985 15240 12019
rect 15182 11951 15240 11985
rect 15182 11917 15194 11951
rect 15228 11917 15240 11951
rect 15182 11883 15240 11917
rect 15182 11849 15194 11883
rect 15228 11849 15240 11883
rect 15182 11815 15240 11849
rect 15182 11781 15194 11815
rect 15228 11781 15240 11815
rect 15182 11747 15240 11781
rect 15182 11713 15194 11747
rect 15228 11713 15240 11747
rect 15182 11679 15240 11713
rect 15182 11645 15194 11679
rect 15228 11645 15240 11679
rect 15182 11611 15240 11645
rect 15182 11577 15194 11611
rect 15228 11577 15240 11611
rect 15182 11543 15240 11577
rect 15182 11509 15194 11543
rect 15228 11509 15240 11543
rect 15182 11475 15240 11509
rect 15182 11441 15194 11475
rect 15228 11441 15240 11475
rect 15182 11407 15240 11441
rect 15182 11373 15194 11407
rect 15228 11373 15240 11407
rect 15182 11339 15240 11373
rect 15182 11305 15194 11339
rect 15228 11305 15240 11339
rect 15182 11271 15240 11305
rect 15182 11237 15194 11271
rect 15228 11237 15240 11271
rect 15182 11203 15240 11237
rect 15182 11169 15194 11203
rect 15228 11169 15240 11203
rect 15182 11135 15240 11169
rect 15182 11101 15194 11135
rect 15228 11101 15240 11135
rect 15182 11070 15240 11101
rect 15270 13039 15328 13070
rect 15270 13005 15282 13039
rect 15316 13005 15328 13039
rect 15270 12971 15328 13005
rect 15270 12937 15282 12971
rect 15316 12937 15328 12971
rect 15270 12903 15328 12937
rect 15270 12869 15282 12903
rect 15316 12869 15328 12903
rect 15270 12835 15328 12869
rect 15270 12801 15282 12835
rect 15316 12801 15328 12835
rect 15270 12767 15328 12801
rect 15270 12733 15282 12767
rect 15316 12733 15328 12767
rect 15270 12699 15328 12733
rect 15270 12665 15282 12699
rect 15316 12665 15328 12699
rect 15270 12631 15328 12665
rect 15270 12597 15282 12631
rect 15316 12597 15328 12631
rect 15270 12563 15328 12597
rect 15270 12529 15282 12563
rect 15316 12529 15328 12563
rect 15270 12495 15328 12529
rect 15270 12461 15282 12495
rect 15316 12461 15328 12495
rect 15270 12427 15328 12461
rect 15270 12393 15282 12427
rect 15316 12393 15328 12427
rect 15270 12359 15328 12393
rect 15270 12325 15282 12359
rect 15316 12325 15328 12359
rect 15270 12291 15328 12325
rect 15270 12257 15282 12291
rect 15316 12257 15328 12291
rect 15270 12223 15328 12257
rect 15270 12189 15282 12223
rect 15316 12189 15328 12223
rect 15270 12155 15328 12189
rect 15270 12121 15282 12155
rect 15316 12121 15328 12155
rect 15270 12087 15328 12121
rect 15270 12053 15282 12087
rect 15316 12053 15328 12087
rect 15270 12019 15328 12053
rect 15270 11985 15282 12019
rect 15316 11985 15328 12019
rect 15270 11951 15328 11985
rect 15270 11917 15282 11951
rect 15316 11917 15328 11951
rect 15270 11883 15328 11917
rect 15270 11849 15282 11883
rect 15316 11849 15328 11883
rect 15270 11815 15328 11849
rect 15270 11781 15282 11815
rect 15316 11781 15328 11815
rect 15270 11747 15328 11781
rect 15270 11713 15282 11747
rect 15316 11713 15328 11747
rect 15270 11679 15328 11713
rect 15270 11645 15282 11679
rect 15316 11645 15328 11679
rect 15270 11611 15328 11645
rect 15270 11577 15282 11611
rect 15316 11577 15328 11611
rect 15270 11543 15328 11577
rect 15270 11509 15282 11543
rect 15316 11509 15328 11543
rect 15270 11475 15328 11509
rect 15270 11441 15282 11475
rect 15316 11441 15328 11475
rect 15270 11407 15328 11441
rect 15270 11373 15282 11407
rect 15316 11373 15328 11407
rect 15270 11339 15328 11373
rect 15270 11305 15282 11339
rect 15316 11305 15328 11339
rect 15270 11271 15328 11305
rect 15270 11237 15282 11271
rect 15316 11237 15328 11271
rect 15270 11203 15328 11237
rect 15270 11169 15282 11203
rect 15316 11169 15328 11203
rect 15270 11135 15328 11169
rect 15270 11101 15282 11135
rect 15316 11101 15328 11135
rect 15270 11070 15328 11101
rect 15358 13039 15416 13070
rect 15358 13005 15370 13039
rect 15404 13005 15416 13039
rect 15358 12971 15416 13005
rect 15358 12937 15370 12971
rect 15404 12937 15416 12971
rect 15358 12903 15416 12937
rect 15358 12869 15370 12903
rect 15404 12869 15416 12903
rect 15358 12835 15416 12869
rect 15358 12801 15370 12835
rect 15404 12801 15416 12835
rect 15358 12767 15416 12801
rect 15358 12733 15370 12767
rect 15404 12733 15416 12767
rect 15358 12699 15416 12733
rect 15358 12665 15370 12699
rect 15404 12665 15416 12699
rect 15358 12631 15416 12665
rect 15358 12597 15370 12631
rect 15404 12597 15416 12631
rect 15358 12563 15416 12597
rect 15358 12529 15370 12563
rect 15404 12529 15416 12563
rect 15358 12495 15416 12529
rect 15358 12461 15370 12495
rect 15404 12461 15416 12495
rect 15358 12427 15416 12461
rect 15358 12393 15370 12427
rect 15404 12393 15416 12427
rect 15358 12359 15416 12393
rect 15358 12325 15370 12359
rect 15404 12325 15416 12359
rect 15358 12291 15416 12325
rect 15358 12257 15370 12291
rect 15404 12257 15416 12291
rect 15358 12223 15416 12257
rect 15358 12189 15370 12223
rect 15404 12189 15416 12223
rect 15358 12155 15416 12189
rect 15358 12121 15370 12155
rect 15404 12121 15416 12155
rect 15358 12087 15416 12121
rect 15358 12053 15370 12087
rect 15404 12053 15416 12087
rect 15358 12019 15416 12053
rect 15358 11985 15370 12019
rect 15404 11985 15416 12019
rect 15358 11951 15416 11985
rect 15358 11917 15370 11951
rect 15404 11917 15416 11951
rect 15358 11883 15416 11917
rect 15358 11849 15370 11883
rect 15404 11849 15416 11883
rect 15358 11815 15416 11849
rect 15358 11781 15370 11815
rect 15404 11781 15416 11815
rect 15358 11747 15416 11781
rect 15358 11713 15370 11747
rect 15404 11713 15416 11747
rect 15358 11679 15416 11713
rect 15358 11645 15370 11679
rect 15404 11645 15416 11679
rect 15358 11611 15416 11645
rect 15358 11577 15370 11611
rect 15404 11577 15416 11611
rect 15358 11543 15416 11577
rect 15358 11509 15370 11543
rect 15404 11509 15416 11543
rect 15358 11475 15416 11509
rect 15358 11441 15370 11475
rect 15404 11441 15416 11475
rect 15358 11407 15416 11441
rect 15358 11373 15370 11407
rect 15404 11373 15416 11407
rect 15358 11339 15416 11373
rect 15358 11305 15370 11339
rect 15404 11305 15416 11339
rect 15358 11271 15416 11305
rect 15358 11237 15370 11271
rect 15404 11237 15416 11271
rect 15358 11203 15416 11237
rect 15358 11169 15370 11203
rect 15404 11169 15416 11203
rect 15358 11135 15416 11169
rect 15358 11101 15370 11135
rect 15404 11101 15416 11135
rect 15358 11070 15416 11101
rect 15446 13039 15504 13070
rect 15446 13005 15458 13039
rect 15492 13005 15504 13039
rect 15446 12971 15504 13005
rect 15446 12937 15458 12971
rect 15492 12937 15504 12971
rect 15446 12903 15504 12937
rect 15446 12869 15458 12903
rect 15492 12869 15504 12903
rect 15446 12835 15504 12869
rect 15446 12801 15458 12835
rect 15492 12801 15504 12835
rect 15446 12767 15504 12801
rect 15446 12733 15458 12767
rect 15492 12733 15504 12767
rect 15446 12699 15504 12733
rect 15446 12665 15458 12699
rect 15492 12665 15504 12699
rect 15446 12631 15504 12665
rect 15446 12597 15458 12631
rect 15492 12597 15504 12631
rect 15446 12563 15504 12597
rect 15446 12529 15458 12563
rect 15492 12529 15504 12563
rect 15446 12495 15504 12529
rect 15446 12461 15458 12495
rect 15492 12461 15504 12495
rect 15446 12427 15504 12461
rect 15446 12393 15458 12427
rect 15492 12393 15504 12427
rect 15446 12359 15504 12393
rect 15446 12325 15458 12359
rect 15492 12325 15504 12359
rect 15446 12291 15504 12325
rect 15446 12257 15458 12291
rect 15492 12257 15504 12291
rect 15446 12223 15504 12257
rect 15446 12189 15458 12223
rect 15492 12189 15504 12223
rect 15446 12155 15504 12189
rect 15446 12121 15458 12155
rect 15492 12121 15504 12155
rect 15446 12087 15504 12121
rect 15446 12053 15458 12087
rect 15492 12053 15504 12087
rect 15446 12019 15504 12053
rect 15446 11985 15458 12019
rect 15492 11985 15504 12019
rect 15446 11951 15504 11985
rect 15446 11917 15458 11951
rect 15492 11917 15504 11951
rect 15446 11883 15504 11917
rect 15446 11849 15458 11883
rect 15492 11849 15504 11883
rect 15446 11815 15504 11849
rect 15446 11781 15458 11815
rect 15492 11781 15504 11815
rect 15446 11747 15504 11781
rect 15446 11713 15458 11747
rect 15492 11713 15504 11747
rect 15446 11679 15504 11713
rect 15446 11645 15458 11679
rect 15492 11645 15504 11679
rect 15446 11611 15504 11645
rect 15446 11577 15458 11611
rect 15492 11577 15504 11611
rect 15446 11543 15504 11577
rect 15446 11509 15458 11543
rect 15492 11509 15504 11543
rect 15446 11475 15504 11509
rect 15446 11441 15458 11475
rect 15492 11441 15504 11475
rect 15446 11407 15504 11441
rect 15446 11373 15458 11407
rect 15492 11373 15504 11407
rect 15446 11339 15504 11373
rect 15446 11305 15458 11339
rect 15492 11305 15504 11339
rect 15446 11271 15504 11305
rect 15446 11237 15458 11271
rect 15492 11237 15504 11271
rect 15446 11203 15504 11237
rect 15446 11169 15458 11203
rect 15492 11169 15504 11203
rect 15446 11135 15504 11169
rect 15446 11101 15458 11135
rect 15492 11101 15504 11135
rect 15446 11070 15504 11101
rect 15534 13039 15592 13070
rect 15534 13005 15546 13039
rect 15580 13005 15592 13039
rect 15534 12971 15592 13005
rect 15534 12937 15546 12971
rect 15580 12937 15592 12971
rect 15534 12903 15592 12937
rect 15534 12869 15546 12903
rect 15580 12869 15592 12903
rect 15534 12835 15592 12869
rect 15534 12801 15546 12835
rect 15580 12801 15592 12835
rect 15534 12767 15592 12801
rect 15534 12733 15546 12767
rect 15580 12733 15592 12767
rect 15534 12699 15592 12733
rect 15534 12665 15546 12699
rect 15580 12665 15592 12699
rect 15534 12631 15592 12665
rect 15534 12597 15546 12631
rect 15580 12597 15592 12631
rect 15534 12563 15592 12597
rect 15534 12529 15546 12563
rect 15580 12529 15592 12563
rect 15534 12495 15592 12529
rect 15534 12461 15546 12495
rect 15580 12461 15592 12495
rect 15534 12427 15592 12461
rect 15534 12393 15546 12427
rect 15580 12393 15592 12427
rect 15534 12359 15592 12393
rect 15534 12325 15546 12359
rect 15580 12325 15592 12359
rect 15534 12291 15592 12325
rect 15534 12257 15546 12291
rect 15580 12257 15592 12291
rect 15534 12223 15592 12257
rect 15534 12189 15546 12223
rect 15580 12189 15592 12223
rect 15534 12155 15592 12189
rect 15534 12121 15546 12155
rect 15580 12121 15592 12155
rect 15534 12087 15592 12121
rect 15534 12053 15546 12087
rect 15580 12053 15592 12087
rect 15534 12019 15592 12053
rect 15534 11985 15546 12019
rect 15580 11985 15592 12019
rect 15534 11951 15592 11985
rect 15534 11917 15546 11951
rect 15580 11917 15592 11951
rect 15534 11883 15592 11917
rect 15534 11849 15546 11883
rect 15580 11849 15592 11883
rect 15534 11815 15592 11849
rect 15534 11781 15546 11815
rect 15580 11781 15592 11815
rect 15534 11747 15592 11781
rect 15534 11713 15546 11747
rect 15580 11713 15592 11747
rect 15534 11679 15592 11713
rect 15534 11645 15546 11679
rect 15580 11645 15592 11679
rect 15534 11611 15592 11645
rect 15534 11577 15546 11611
rect 15580 11577 15592 11611
rect 15534 11543 15592 11577
rect 15534 11509 15546 11543
rect 15580 11509 15592 11543
rect 15534 11475 15592 11509
rect 15534 11441 15546 11475
rect 15580 11441 15592 11475
rect 15534 11407 15592 11441
rect 15534 11373 15546 11407
rect 15580 11373 15592 11407
rect 15534 11339 15592 11373
rect 15534 11305 15546 11339
rect 15580 11305 15592 11339
rect 15534 11271 15592 11305
rect 15534 11237 15546 11271
rect 15580 11237 15592 11271
rect 15534 11203 15592 11237
rect 15534 11169 15546 11203
rect 15580 11169 15592 11203
rect 15534 11135 15592 11169
rect 15534 11101 15546 11135
rect 15580 11101 15592 11135
rect 15534 11070 15592 11101
rect 15622 13039 15680 13070
rect 15622 13005 15634 13039
rect 15668 13005 15680 13039
rect 15622 12971 15680 13005
rect 15622 12937 15634 12971
rect 15668 12937 15680 12971
rect 15622 12903 15680 12937
rect 15622 12869 15634 12903
rect 15668 12869 15680 12903
rect 15622 12835 15680 12869
rect 15622 12801 15634 12835
rect 15668 12801 15680 12835
rect 15622 12767 15680 12801
rect 15622 12733 15634 12767
rect 15668 12733 15680 12767
rect 15622 12699 15680 12733
rect 15622 12665 15634 12699
rect 15668 12665 15680 12699
rect 15622 12631 15680 12665
rect 15622 12597 15634 12631
rect 15668 12597 15680 12631
rect 15622 12563 15680 12597
rect 15622 12529 15634 12563
rect 15668 12529 15680 12563
rect 15622 12495 15680 12529
rect 15622 12461 15634 12495
rect 15668 12461 15680 12495
rect 15622 12427 15680 12461
rect 15622 12393 15634 12427
rect 15668 12393 15680 12427
rect 15622 12359 15680 12393
rect 15622 12325 15634 12359
rect 15668 12325 15680 12359
rect 15622 12291 15680 12325
rect 15622 12257 15634 12291
rect 15668 12257 15680 12291
rect 15622 12223 15680 12257
rect 15622 12189 15634 12223
rect 15668 12189 15680 12223
rect 15622 12155 15680 12189
rect 15622 12121 15634 12155
rect 15668 12121 15680 12155
rect 15622 12087 15680 12121
rect 15622 12053 15634 12087
rect 15668 12053 15680 12087
rect 15622 12019 15680 12053
rect 15622 11985 15634 12019
rect 15668 11985 15680 12019
rect 15622 11951 15680 11985
rect 15622 11917 15634 11951
rect 15668 11917 15680 11951
rect 15622 11883 15680 11917
rect 15622 11849 15634 11883
rect 15668 11849 15680 11883
rect 15622 11815 15680 11849
rect 15622 11781 15634 11815
rect 15668 11781 15680 11815
rect 15622 11747 15680 11781
rect 15622 11713 15634 11747
rect 15668 11713 15680 11747
rect 15622 11679 15680 11713
rect 15622 11645 15634 11679
rect 15668 11645 15680 11679
rect 15622 11611 15680 11645
rect 15622 11577 15634 11611
rect 15668 11577 15680 11611
rect 15622 11543 15680 11577
rect 15622 11509 15634 11543
rect 15668 11509 15680 11543
rect 15622 11475 15680 11509
rect 15622 11441 15634 11475
rect 15668 11441 15680 11475
rect 15622 11407 15680 11441
rect 15622 11373 15634 11407
rect 15668 11373 15680 11407
rect 15622 11339 15680 11373
rect 15622 11305 15634 11339
rect 15668 11305 15680 11339
rect 15622 11271 15680 11305
rect 15622 11237 15634 11271
rect 15668 11237 15680 11271
rect 15622 11203 15680 11237
rect 15622 11169 15634 11203
rect 15668 11169 15680 11203
rect 15622 11135 15680 11169
rect 15622 11101 15634 11135
rect 15668 11101 15680 11135
rect 15622 11070 15680 11101
rect 15710 13039 15768 13070
rect 15710 13005 15722 13039
rect 15756 13005 15768 13039
rect 15710 12971 15768 13005
rect 15710 12937 15722 12971
rect 15756 12937 15768 12971
rect 15710 12903 15768 12937
rect 15710 12869 15722 12903
rect 15756 12869 15768 12903
rect 15710 12835 15768 12869
rect 15710 12801 15722 12835
rect 15756 12801 15768 12835
rect 15710 12767 15768 12801
rect 15710 12733 15722 12767
rect 15756 12733 15768 12767
rect 15710 12699 15768 12733
rect 15710 12665 15722 12699
rect 15756 12665 15768 12699
rect 15710 12631 15768 12665
rect 15710 12597 15722 12631
rect 15756 12597 15768 12631
rect 15710 12563 15768 12597
rect 15710 12529 15722 12563
rect 15756 12529 15768 12563
rect 15710 12495 15768 12529
rect 15710 12461 15722 12495
rect 15756 12461 15768 12495
rect 15710 12427 15768 12461
rect 15710 12393 15722 12427
rect 15756 12393 15768 12427
rect 15710 12359 15768 12393
rect 15710 12325 15722 12359
rect 15756 12325 15768 12359
rect 15710 12291 15768 12325
rect 15710 12257 15722 12291
rect 15756 12257 15768 12291
rect 15710 12223 15768 12257
rect 15710 12189 15722 12223
rect 15756 12189 15768 12223
rect 15710 12155 15768 12189
rect 15710 12121 15722 12155
rect 15756 12121 15768 12155
rect 15710 12087 15768 12121
rect 15710 12053 15722 12087
rect 15756 12053 15768 12087
rect 15710 12019 15768 12053
rect 15710 11985 15722 12019
rect 15756 11985 15768 12019
rect 15710 11951 15768 11985
rect 15710 11917 15722 11951
rect 15756 11917 15768 11951
rect 15710 11883 15768 11917
rect 15710 11849 15722 11883
rect 15756 11849 15768 11883
rect 15710 11815 15768 11849
rect 15710 11781 15722 11815
rect 15756 11781 15768 11815
rect 15710 11747 15768 11781
rect 15710 11713 15722 11747
rect 15756 11713 15768 11747
rect 15710 11679 15768 11713
rect 15710 11645 15722 11679
rect 15756 11645 15768 11679
rect 15710 11611 15768 11645
rect 15710 11577 15722 11611
rect 15756 11577 15768 11611
rect 15710 11543 15768 11577
rect 15710 11509 15722 11543
rect 15756 11509 15768 11543
rect 15710 11475 15768 11509
rect 15710 11441 15722 11475
rect 15756 11441 15768 11475
rect 15710 11407 15768 11441
rect 15710 11373 15722 11407
rect 15756 11373 15768 11407
rect 15710 11339 15768 11373
rect 15710 11305 15722 11339
rect 15756 11305 15768 11339
rect 15710 11271 15768 11305
rect 15710 11237 15722 11271
rect 15756 11237 15768 11271
rect 15710 11203 15768 11237
rect 15710 11169 15722 11203
rect 15756 11169 15768 11203
rect 15710 11135 15768 11169
rect 15710 11101 15722 11135
rect 15756 11101 15768 11135
rect 15710 11070 15768 11101
rect 15798 13039 15856 13070
rect 15798 13005 15810 13039
rect 15844 13005 15856 13039
rect 15798 12971 15856 13005
rect 15798 12937 15810 12971
rect 15844 12937 15856 12971
rect 15798 12903 15856 12937
rect 15798 12869 15810 12903
rect 15844 12869 15856 12903
rect 15798 12835 15856 12869
rect 15798 12801 15810 12835
rect 15844 12801 15856 12835
rect 15798 12767 15856 12801
rect 15798 12733 15810 12767
rect 15844 12733 15856 12767
rect 15798 12699 15856 12733
rect 15798 12665 15810 12699
rect 15844 12665 15856 12699
rect 15798 12631 15856 12665
rect 15798 12597 15810 12631
rect 15844 12597 15856 12631
rect 15798 12563 15856 12597
rect 15798 12529 15810 12563
rect 15844 12529 15856 12563
rect 15798 12495 15856 12529
rect 15798 12461 15810 12495
rect 15844 12461 15856 12495
rect 15798 12427 15856 12461
rect 15798 12393 15810 12427
rect 15844 12393 15856 12427
rect 15798 12359 15856 12393
rect 15798 12325 15810 12359
rect 15844 12325 15856 12359
rect 15798 12291 15856 12325
rect 15798 12257 15810 12291
rect 15844 12257 15856 12291
rect 15798 12223 15856 12257
rect 15798 12189 15810 12223
rect 15844 12189 15856 12223
rect 15798 12155 15856 12189
rect 15798 12121 15810 12155
rect 15844 12121 15856 12155
rect 15798 12087 15856 12121
rect 15798 12053 15810 12087
rect 15844 12053 15856 12087
rect 15798 12019 15856 12053
rect 15798 11985 15810 12019
rect 15844 11985 15856 12019
rect 15798 11951 15856 11985
rect 15798 11917 15810 11951
rect 15844 11917 15856 11951
rect 15798 11883 15856 11917
rect 15798 11849 15810 11883
rect 15844 11849 15856 11883
rect 15798 11815 15856 11849
rect 15798 11781 15810 11815
rect 15844 11781 15856 11815
rect 15798 11747 15856 11781
rect 15798 11713 15810 11747
rect 15844 11713 15856 11747
rect 15798 11679 15856 11713
rect 15798 11645 15810 11679
rect 15844 11645 15856 11679
rect 15798 11611 15856 11645
rect 15798 11577 15810 11611
rect 15844 11577 15856 11611
rect 15798 11543 15856 11577
rect 15798 11509 15810 11543
rect 15844 11509 15856 11543
rect 15798 11475 15856 11509
rect 15798 11441 15810 11475
rect 15844 11441 15856 11475
rect 15798 11407 15856 11441
rect 15798 11373 15810 11407
rect 15844 11373 15856 11407
rect 15798 11339 15856 11373
rect 15798 11305 15810 11339
rect 15844 11305 15856 11339
rect 15798 11271 15856 11305
rect 15798 11237 15810 11271
rect 15844 11237 15856 11271
rect 15798 11203 15856 11237
rect 15798 11169 15810 11203
rect 15844 11169 15856 11203
rect 15798 11135 15856 11169
rect 15798 11101 15810 11135
rect 15844 11101 15856 11135
rect 15798 11070 15856 11101
rect 15886 13039 15944 13070
rect 15886 13005 15898 13039
rect 15932 13005 15944 13039
rect 15886 12971 15944 13005
rect 15886 12937 15898 12971
rect 15932 12937 15944 12971
rect 15886 12903 15944 12937
rect 15886 12869 15898 12903
rect 15932 12869 15944 12903
rect 15886 12835 15944 12869
rect 15886 12801 15898 12835
rect 15932 12801 15944 12835
rect 15886 12767 15944 12801
rect 15886 12733 15898 12767
rect 15932 12733 15944 12767
rect 15886 12699 15944 12733
rect 15886 12665 15898 12699
rect 15932 12665 15944 12699
rect 15886 12631 15944 12665
rect 15886 12597 15898 12631
rect 15932 12597 15944 12631
rect 15886 12563 15944 12597
rect 15886 12529 15898 12563
rect 15932 12529 15944 12563
rect 15886 12495 15944 12529
rect 15886 12461 15898 12495
rect 15932 12461 15944 12495
rect 15886 12427 15944 12461
rect 15886 12393 15898 12427
rect 15932 12393 15944 12427
rect 15886 12359 15944 12393
rect 15886 12325 15898 12359
rect 15932 12325 15944 12359
rect 15886 12291 15944 12325
rect 15886 12257 15898 12291
rect 15932 12257 15944 12291
rect 15886 12223 15944 12257
rect 15886 12189 15898 12223
rect 15932 12189 15944 12223
rect 15886 12155 15944 12189
rect 15886 12121 15898 12155
rect 15932 12121 15944 12155
rect 15886 12087 15944 12121
rect 15886 12053 15898 12087
rect 15932 12053 15944 12087
rect 15886 12019 15944 12053
rect 15886 11985 15898 12019
rect 15932 11985 15944 12019
rect 15886 11951 15944 11985
rect 15886 11917 15898 11951
rect 15932 11917 15944 11951
rect 15886 11883 15944 11917
rect 15886 11849 15898 11883
rect 15932 11849 15944 11883
rect 15886 11815 15944 11849
rect 15886 11781 15898 11815
rect 15932 11781 15944 11815
rect 15886 11747 15944 11781
rect 15886 11713 15898 11747
rect 15932 11713 15944 11747
rect 15886 11679 15944 11713
rect 15886 11645 15898 11679
rect 15932 11645 15944 11679
rect 15886 11611 15944 11645
rect 15886 11577 15898 11611
rect 15932 11577 15944 11611
rect 15886 11543 15944 11577
rect 15886 11509 15898 11543
rect 15932 11509 15944 11543
rect 15886 11475 15944 11509
rect 15886 11441 15898 11475
rect 15932 11441 15944 11475
rect 15886 11407 15944 11441
rect 15886 11373 15898 11407
rect 15932 11373 15944 11407
rect 15886 11339 15944 11373
rect 15886 11305 15898 11339
rect 15932 11305 15944 11339
rect 15886 11271 15944 11305
rect 15886 11237 15898 11271
rect 15932 11237 15944 11271
rect 15886 11203 15944 11237
rect 15886 11169 15898 11203
rect 15932 11169 15944 11203
rect 15886 11135 15944 11169
rect 15886 11101 15898 11135
rect 15932 11101 15944 11135
rect 15886 11070 15944 11101
rect 15974 13039 16032 13070
rect 15974 13005 15986 13039
rect 16020 13005 16032 13039
rect 15974 12971 16032 13005
rect 15974 12937 15986 12971
rect 16020 12937 16032 12971
rect 15974 12903 16032 12937
rect 15974 12869 15986 12903
rect 16020 12869 16032 12903
rect 15974 12835 16032 12869
rect 15974 12801 15986 12835
rect 16020 12801 16032 12835
rect 15974 12767 16032 12801
rect 15974 12733 15986 12767
rect 16020 12733 16032 12767
rect 15974 12699 16032 12733
rect 15974 12665 15986 12699
rect 16020 12665 16032 12699
rect 15974 12631 16032 12665
rect 15974 12597 15986 12631
rect 16020 12597 16032 12631
rect 15974 12563 16032 12597
rect 15974 12529 15986 12563
rect 16020 12529 16032 12563
rect 15974 12495 16032 12529
rect 15974 12461 15986 12495
rect 16020 12461 16032 12495
rect 15974 12427 16032 12461
rect 15974 12393 15986 12427
rect 16020 12393 16032 12427
rect 15974 12359 16032 12393
rect 15974 12325 15986 12359
rect 16020 12325 16032 12359
rect 15974 12291 16032 12325
rect 15974 12257 15986 12291
rect 16020 12257 16032 12291
rect 15974 12223 16032 12257
rect 15974 12189 15986 12223
rect 16020 12189 16032 12223
rect 15974 12155 16032 12189
rect 15974 12121 15986 12155
rect 16020 12121 16032 12155
rect 15974 12087 16032 12121
rect 15974 12053 15986 12087
rect 16020 12053 16032 12087
rect 15974 12019 16032 12053
rect 15974 11985 15986 12019
rect 16020 11985 16032 12019
rect 15974 11951 16032 11985
rect 15974 11917 15986 11951
rect 16020 11917 16032 11951
rect 15974 11883 16032 11917
rect 15974 11849 15986 11883
rect 16020 11849 16032 11883
rect 15974 11815 16032 11849
rect 15974 11781 15986 11815
rect 16020 11781 16032 11815
rect 15974 11747 16032 11781
rect 15974 11713 15986 11747
rect 16020 11713 16032 11747
rect 15974 11679 16032 11713
rect 15974 11645 15986 11679
rect 16020 11645 16032 11679
rect 15974 11611 16032 11645
rect 15974 11577 15986 11611
rect 16020 11577 16032 11611
rect 15974 11543 16032 11577
rect 15974 11509 15986 11543
rect 16020 11509 16032 11543
rect 15974 11475 16032 11509
rect 15974 11441 15986 11475
rect 16020 11441 16032 11475
rect 15974 11407 16032 11441
rect 15974 11373 15986 11407
rect 16020 11373 16032 11407
rect 15974 11339 16032 11373
rect 15974 11305 15986 11339
rect 16020 11305 16032 11339
rect 15974 11271 16032 11305
rect 15974 11237 15986 11271
rect 16020 11237 16032 11271
rect 15974 11203 16032 11237
rect 15974 11169 15986 11203
rect 16020 11169 16032 11203
rect 15974 11135 16032 11169
rect 15974 11101 15986 11135
rect 16020 11101 16032 11135
rect 15974 11070 16032 11101
rect 16062 13039 16120 13070
rect 16062 13005 16074 13039
rect 16108 13005 16120 13039
rect 16062 12971 16120 13005
rect 16062 12937 16074 12971
rect 16108 12937 16120 12971
rect 16062 12903 16120 12937
rect 16062 12869 16074 12903
rect 16108 12869 16120 12903
rect 16062 12835 16120 12869
rect 16062 12801 16074 12835
rect 16108 12801 16120 12835
rect 16062 12767 16120 12801
rect 16062 12733 16074 12767
rect 16108 12733 16120 12767
rect 16062 12699 16120 12733
rect 16062 12665 16074 12699
rect 16108 12665 16120 12699
rect 16062 12631 16120 12665
rect 16062 12597 16074 12631
rect 16108 12597 16120 12631
rect 16062 12563 16120 12597
rect 16062 12529 16074 12563
rect 16108 12529 16120 12563
rect 16062 12495 16120 12529
rect 16062 12461 16074 12495
rect 16108 12461 16120 12495
rect 16062 12427 16120 12461
rect 16062 12393 16074 12427
rect 16108 12393 16120 12427
rect 16062 12359 16120 12393
rect 16062 12325 16074 12359
rect 16108 12325 16120 12359
rect 16062 12291 16120 12325
rect 16062 12257 16074 12291
rect 16108 12257 16120 12291
rect 16062 12223 16120 12257
rect 16062 12189 16074 12223
rect 16108 12189 16120 12223
rect 16062 12155 16120 12189
rect 16062 12121 16074 12155
rect 16108 12121 16120 12155
rect 16062 12087 16120 12121
rect 16062 12053 16074 12087
rect 16108 12053 16120 12087
rect 16062 12019 16120 12053
rect 16062 11985 16074 12019
rect 16108 11985 16120 12019
rect 16062 11951 16120 11985
rect 16062 11917 16074 11951
rect 16108 11917 16120 11951
rect 16062 11883 16120 11917
rect 16062 11849 16074 11883
rect 16108 11849 16120 11883
rect 16062 11815 16120 11849
rect 16062 11781 16074 11815
rect 16108 11781 16120 11815
rect 16062 11747 16120 11781
rect 16062 11713 16074 11747
rect 16108 11713 16120 11747
rect 16062 11679 16120 11713
rect 16062 11645 16074 11679
rect 16108 11645 16120 11679
rect 16062 11611 16120 11645
rect 16062 11577 16074 11611
rect 16108 11577 16120 11611
rect 16062 11543 16120 11577
rect 16062 11509 16074 11543
rect 16108 11509 16120 11543
rect 16062 11475 16120 11509
rect 16062 11441 16074 11475
rect 16108 11441 16120 11475
rect 16062 11407 16120 11441
rect 16062 11373 16074 11407
rect 16108 11373 16120 11407
rect 16062 11339 16120 11373
rect 16062 11305 16074 11339
rect 16108 11305 16120 11339
rect 16062 11271 16120 11305
rect 16062 11237 16074 11271
rect 16108 11237 16120 11271
rect 16062 11203 16120 11237
rect 16062 11169 16074 11203
rect 16108 11169 16120 11203
rect 16062 11135 16120 11169
rect 16062 11101 16074 11135
rect 16108 11101 16120 11135
rect 16062 11070 16120 11101
rect 16150 13039 16208 13070
rect 16150 13005 16162 13039
rect 16196 13005 16208 13039
rect 16150 12971 16208 13005
rect 16150 12937 16162 12971
rect 16196 12937 16208 12971
rect 16150 12903 16208 12937
rect 16150 12869 16162 12903
rect 16196 12869 16208 12903
rect 16150 12835 16208 12869
rect 16150 12801 16162 12835
rect 16196 12801 16208 12835
rect 16150 12767 16208 12801
rect 16150 12733 16162 12767
rect 16196 12733 16208 12767
rect 16150 12699 16208 12733
rect 16150 12665 16162 12699
rect 16196 12665 16208 12699
rect 16150 12631 16208 12665
rect 16150 12597 16162 12631
rect 16196 12597 16208 12631
rect 16150 12563 16208 12597
rect 16150 12529 16162 12563
rect 16196 12529 16208 12563
rect 16150 12495 16208 12529
rect 16150 12461 16162 12495
rect 16196 12461 16208 12495
rect 16150 12427 16208 12461
rect 16150 12393 16162 12427
rect 16196 12393 16208 12427
rect 16150 12359 16208 12393
rect 16150 12325 16162 12359
rect 16196 12325 16208 12359
rect 16150 12291 16208 12325
rect 16150 12257 16162 12291
rect 16196 12257 16208 12291
rect 16150 12223 16208 12257
rect 16150 12189 16162 12223
rect 16196 12189 16208 12223
rect 16150 12155 16208 12189
rect 16150 12121 16162 12155
rect 16196 12121 16208 12155
rect 16150 12087 16208 12121
rect 16150 12053 16162 12087
rect 16196 12053 16208 12087
rect 16150 12019 16208 12053
rect 16150 11985 16162 12019
rect 16196 11985 16208 12019
rect 16150 11951 16208 11985
rect 16150 11917 16162 11951
rect 16196 11917 16208 11951
rect 16150 11883 16208 11917
rect 16150 11849 16162 11883
rect 16196 11849 16208 11883
rect 16150 11815 16208 11849
rect 16150 11781 16162 11815
rect 16196 11781 16208 11815
rect 16150 11747 16208 11781
rect 16150 11713 16162 11747
rect 16196 11713 16208 11747
rect 16150 11679 16208 11713
rect 16150 11645 16162 11679
rect 16196 11645 16208 11679
rect 16150 11611 16208 11645
rect 16150 11577 16162 11611
rect 16196 11577 16208 11611
rect 16150 11543 16208 11577
rect 16150 11509 16162 11543
rect 16196 11509 16208 11543
rect 16150 11475 16208 11509
rect 16150 11441 16162 11475
rect 16196 11441 16208 11475
rect 16150 11407 16208 11441
rect 16150 11373 16162 11407
rect 16196 11373 16208 11407
rect 16150 11339 16208 11373
rect 16150 11305 16162 11339
rect 16196 11305 16208 11339
rect 16150 11271 16208 11305
rect 16150 11237 16162 11271
rect 16196 11237 16208 11271
rect 16150 11203 16208 11237
rect 16150 11169 16162 11203
rect 16196 11169 16208 11203
rect 16150 11135 16208 11169
rect 16150 11101 16162 11135
rect 16196 11101 16208 11135
rect 16150 11070 16208 11101
rect 16238 13039 16296 13070
rect 16238 13005 16250 13039
rect 16284 13005 16296 13039
rect 16238 12971 16296 13005
rect 16238 12937 16250 12971
rect 16284 12937 16296 12971
rect 16238 12903 16296 12937
rect 16238 12869 16250 12903
rect 16284 12869 16296 12903
rect 16238 12835 16296 12869
rect 16238 12801 16250 12835
rect 16284 12801 16296 12835
rect 16238 12767 16296 12801
rect 16238 12733 16250 12767
rect 16284 12733 16296 12767
rect 16238 12699 16296 12733
rect 16238 12665 16250 12699
rect 16284 12665 16296 12699
rect 16238 12631 16296 12665
rect 16238 12597 16250 12631
rect 16284 12597 16296 12631
rect 16238 12563 16296 12597
rect 16238 12529 16250 12563
rect 16284 12529 16296 12563
rect 16238 12495 16296 12529
rect 16238 12461 16250 12495
rect 16284 12461 16296 12495
rect 16238 12427 16296 12461
rect 16238 12393 16250 12427
rect 16284 12393 16296 12427
rect 16238 12359 16296 12393
rect 16238 12325 16250 12359
rect 16284 12325 16296 12359
rect 16238 12291 16296 12325
rect 16238 12257 16250 12291
rect 16284 12257 16296 12291
rect 16238 12223 16296 12257
rect 16238 12189 16250 12223
rect 16284 12189 16296 12223
rect 16238 12155 16296 12189
rect 16238 12121 16250 12155
rect 16284 12121 16296 12155
rect 16238 12087 16296 12121
rect 16238 12053 16250 12087
rect 16284 12053 16296 12087
rect 16238 12019 16296 12053
rect 16238 11985 16250 12019
rect 16284 11985 16296 12019
rect 16238 11951 16296 11985
rect 16238 11917 16250 11951
rect 16284 11917 16296 11951
rect 16238 11883 16296 11917
rect 16238 11849 16250 11883
rect 16284 11849 16296 11883
rect 16238 11815 16296 11849
rect 16238 11781 16250 11815
rect 16284 11781 16296 11815
rect 16238 11747 16296 11781
rect 16238 11713 16250 11747
rect 16284 11713 16296 11747
rect 16238 11679 16296 11713
rect 16238 11645 16250 11679
rect 16284 11645 16296 11679
rect 16238 11611 16296 11645
rect 16238 11577 16250 11611
rect 16284 11577 16296 11611
rect 16238 11543 16296 11577
rect 16238 11509 16250 11543
rect 16284 11509 16296 11543
rect 16238 11475 16296 11509
rect 16238 11441 16250 11475
rect 16284 11441 16296 11475
rect 16238 11407 16296 11441
rect 16238 11373 16250 11407
rect 16284 11373 16296 11407
rect 16238 11339 16296 11373
rect 16238 11305 16250 11339
rect 16284 11305 16296 11339
rect 16238 11271 16296 11305
rect 16238 11237 16250 11271
rect 16284 11237 16296 11271
rect 16238 11203 16296 11237
rect 16238 11169 16250 11203
rect 16284 11169 16296 11203
rect 16238 11135 16296 11169
rect 16238 11101 16250 11135
rect 16284 11101 16296 11135
rect 16238 11070 16296 11101
rect 16326 13039 16384 13070
rect 16326 13005 16338 13039
rect 16372 13005 16384 13039
rect 16326 12971 16384 13005
rect 16326 12937 16338 12971
rect 16372 12937 16384 12971
rect 16326 12903 16384 12937
rect 16326 12869 16338 12903
rect 16372 12869 16384 12903
rect 16326 12835 16384 12869
rect 16326 12801 16338 12835
rect 16372 12801 16384 12835
rect 16326 12767 16384 12801
rect 16326 12733 16338 12767
rect 16372 12733 16384 12767
rect 16326 12699 16384 12733
rect 16326 12665 16338 12699
rect 16372 12665 16384 12699
rect 16326 12631 16384 12665
rect 16326 12597 16338 12631
rect 16372 12597 16384 12631
rect 16326 12563 16384 12597
rect 16326 12529 16338 12563
rect 16372 12529 16384 12563
rect 16326 12495 16384 12529
rect 16326 12461 16338 12495
rect 16372 12461 16384 12495
rect 16326 12427 16384 12461
rect 16326 12393 16338 12427
rect 16372 12393 16384 12427
rect 16326 12359 16384 12393
rect 16326 12325 16338 12359
rect 16372 12325 16384 12359
rect 16326 12291 16384 12325
rect 16326 12257 16338 12291
rect 16372 12257 16384 12291
rect 16326 12223 16384 12257
rect 16326 12189 16338 12223
rect 16372 12189 16384 12223
rect 16326 12155 16384 12189
rect 16326 12121 16338 12155
rect 16372 12121 16384 12155
rect 16326 12087 16384 12121
rect 16326 12053 16338 12087
rect 16372 12053 16384 12087
rect 16326 12019 16384 12053
rect 16326 11985 16338 12019
rect 16372 11985 16384 12019
rect 16326 11951 16384 11985
rect 16326 11917 16338 11951
rect 16372 11917 16384 11951
rect 16326 11883 16384 11917
rect 16326 11849 16338 11883
rect 16372 11849 16384 11883
rect 16326 11815 16384 11849
rect 16326 11781 16338 11815
rect 16372 11781 16384 11815
rect 16326 11747 16384 11781
rect 16326 11713 16338 11747
rect 16372 11713 16384 11747
rect 16326 11679 16384 11713
rect 16326 11645 16338 11679
rect 16372 11645 16384 11679
rect 16326 11611 16384 11645
rect 16326 11577 16338 11611
rect 16372 11577 16384 11611
rect 16326 11543 16384 11577
rect 16326 11509 16338 11543
rect 16372 11509 16384 11543
rect 16326 11475 16384 11509
rect 16326 11441 16338 11475
rect 16372 11441 16384 11475
rect 16326 11407 16384 11441
rect 16326 11373 16338 11407
rect 16372 11373 16384 11407
rect 16326 11339 16384 11373
rect 16326 11305 16338 11339
rect 16372 11305 16384 11339
rect 16326 11271 16384 11305
rect 16326 11237 16338 11271
rect 16372 11237 16384 11271
rect 16326 11203 16384 11237
rect 16326 11169 16338 11203
rect 16372 11169 16384 11203
rect 16326 11135 16384 11169
rect 16326 11101 16338 11135
rect 16372 11101 16384 11135
rect 16326 11070 16384 11101
rect 16414 13039 16472 13070
rect 16414 13005 16426 13039
rect 16460 13005 16472 13039
rect 16414 12971 16472 13005
rect 16414 12937 16426 12971
rect 16460 12937 16472 12971
rect 16414 12903 16472 12937
rect 16414 12869 16426 12903
rect 16460 12869 16472 12903
rect 16414 12835 16472 12869
rect 16414 12801 16426 12835
rect 16460 12801 16472 12835
rect 16414 12767 16472 12801
rect 16414 12733 16426 12767
rect 16460 12733 16472 12767
rect 16414 12699 16472 12733
rect 16414 12665 16426 12699
rect 16460 12665 16472 12699
rect 16414 12631 16472 12665
rect 16414 12597 16426 12631
rect 16460 12597 16472 12631
rect 16414 12563 16472 12597
rect 16414 12529 16426 12563
rect 16460 12529 16472 12563
rect 16414 12495 16472 12529
rect 16414 12461 16426 12495
rect 16460 12461 16472 12495
rect 16414 12427 16472 12461
rect 16414 12393 16426 12427
rect 16460 12393 16472 12427
rect 16414 12359 16472 12393
rect 16414 12325 16426 12359
rect 16460 12325 16472 12359
rect 16414 12291 16472 12325
rect 16414 12257 16426 12291
rect 16460 12257 16472 12291
rect 16414 12223 16472 12257
rect 16414 12189 16426 12223
rect 16460 12189 16472 12223
rect 16414 12155 16472 12189
rect 16414 12121 16426 12155
rect 16460 12121 16472 12155
rect 16414 12087 16472 12121
rect 16414 12053 16426 12087
rect 16460 12053 16472 12087
rect 16414 12019 16472 12053
rect 16414 11985 16426 12019
rect 16460 11985 16472 12019
rect 16414 11951 16472 11985
rect 16414 11917 16426 11951
rect 16460 11917 16472 11951
rect 16414 11883 16472 11917
rect 16414 11849 16426 11883
rect 16460 11849 16472 11883
rect 16414 11815 16472 11849
rect 16414 11781 16426 11815
rect 16460 11781 16472 11815
rect 16414 11747 16472 11781
rect 16414 11713 16426 11747
rect 16460 11713 16472 11747
rect 16414 11679 16472 11713
rect 16414 11645 16426 11679
rect 16460 11645 16472 11679
rect 16414 11611 16472 11645
rect 16414 11577 16426 11611
rect 16460 11577 16472 11611
rect 16414 11543 16472 11577
rect 16414 11509 16426 11543
rect 16460 11509 16472 11543
rect 16414 11475 16472 11509
rect 16414 11441 16426 11475
rect 16460 11441 16472 11475
rect 16414 11407 16472 11441
rect 16414 11373 16426 11407
rect 16460 11373 16472 11407
rect 16414 11339 16472 11373
rect 16414 11305 16426 11339
rect 16460 11305 16472 11339
rect 16414 11271 16472 11305
rect 16414 11237 16426 11271
rect 16460 11237 16472 11271
rect 16414 11203 16472 11237
rect 16414 11169 16426 11203
rect 16460 11169 16472 11203
rect 16414 11135 16472 11169
rect 16414 11101 16426 11135
rect 16460 11101 16472 11135
rect 16414 11070 16472 11101
rect 16502 13039 16560 13070
rect 16502 13005 16514 13039
rect 16548 13005 16560 13039
rect 16502 12971 16560 13005
rect 16502 12937 16514 12971
rect 16548 12937 16560 12971
rect 16502 12903 16560 12937
rect 16502 12869 16514 12903
rect 16548 12869 16560 12903
rect 16502 12835 16560 12869
rect 16502 12801 16514 12835
rect 16548 12801 16560 12835
rect 16502 12767 16560 12801
rect 16502 12733 16514 12767
rect 16548 12733 16560 12767
rect 16502 12699 16560 12733
rect 16502 12665 16514 12699
rect 16548 12665 16560 12699
rect 16502 12631 16560 12665
rect 16502 12597 16514 12631
rect 16548 12597 16560 12631
rect 16502 12563 16560 12597
rect 16502 12529 16514 12563
rect 16548 12529 16560 12563
rect 16502 12495 16560 12529
rect 16502 12461 16514 12495
rect 16548 12461 16560 12495
rect 16502 12427 16560 12461
rect 16502 12393 16514 12427
rect 16548 12393 16560 12427
rect 16502 12359 16560 12393
rect 16502 12325 16514 12359
rect 16548 12325 16560 12359
rect 16502 12291 16560 12325
rect 16502 12257 16514 12291
rect 16548 12257 16560 12291
rect 16502 12223 16560 12257
rect 16502 12189 16514 12223
rect 16548 12189 16560 12223
rect 16502 12155 16560 12189
rect 16502 12121 16514 12155
rect 16548 12121 16560 12155
rect 16502 12087 16560 12121
rect 16502 12053 16514 12087
rect 16548 12053 16560 12087
rect 16502 12019 16560 12053
rect 16502 11985 16514 12019
rect 16548 11985 16560 12019
rect 16502 11951 16560 11985
rect 16502 11917 16514 11951
rect 16548 11917 16560 11951
rect 16502 11883 16560 11917
rect 16502 11849 16514 11883
rect 16548 11849 16560 11883
rect 16502 11815 16560 11849
rect 16502 11781 16514 11815
rect 16548 11781 16560 11815
rect 16502 11747 16560 11781
rect 16502 11713 16514 11747
rect 16548 11713 16560 11747
rect 16502 11679 16560 11713
rect 16502 11645 16514 11679
rect 16548 11645 16560 11679
rect 16502 11611 16560 11645
rect 16502 11577 16514 11611
rect 16548 11577 16560 11611
rect 16502 11543 16560 11577
rect 16502 11509 16514 11543
rect 16548 11509 16560 11543
rect 16502 11475 16560 11509
rect 16502 11441 16514 11475
rect 16548 11441 16560 11475
rect 16502 11407 16560 11441
rect 16502 11373 16514 11407
rect 16548 11373 16560 11407
rect 16502 11339 16560 11373
rect 16502 11305 16514 11339
rect 16548 11305 16560 11339
rect 16502 11271 16560 11305
rect 16502 11237 16514 11271
rect 16548 11237 16560 11271
rect 16502 11203 16560 11237
rect 16502 11169 16514 11203
rect 16548 11169 16560 11203
rect 16502 11135 16560 11169
rect 16502 11101 16514 11135
rect 16548 11101 16560 11135
rect 16502 11070 16560 11101
rect 16590 13039 16648 13070
rect 16590 13005 16602 13039
rect 16636 13005 16648 13039
rect 16590 12971 16648 13005
rect 16590 12937 16602 12971
rect 16636 12937 16648 12971
rect 16590 12903 16648 12937
rect 16590 12869 16602 12903
rect 16636 12869 16648 12903
rect 16590 12835 16648 12869
rect 16590 12801 16602 12835
rect 16636 12801 16648 12835
rect 16590 12767 16648 12801
rect 16590 12733 16602 12767
rect 16636 12733 16648 12767
rect 16590 12699 16648 12733
rect 16590 12665 16602 12699
rect 16636 12665 16648 12699
rect 16590 12631 16648 12665
rect 16590 12597 16602 12631
rect 16636 12597 16648 12631
rect 16590 12563 16648 12597
rect 16590 12529 16602 12563
rect 16636 12529 16648 12563
rect 16590 12495 16648 12529
rect 16590 12461 16602 12495
rect 16636 12461 16648 12495
rect 16590 12427 16648 12461
rect 16590 12393 16602 12427
rect 16636 12393 16648 12427
rect 16590 12359 16648 12393
rect 16590 12325 16602 12359
rect 16636 12325 16648 12359
rect 16590 12291 16648 12325
rect 16590 12257 16602 12291
rect 16636 12257 16648 12291
rect 16590 12223 16648 12257
rect 16590 12189 16602 12223
rect 16636 12189 16648 12223
rect 16590 12155 16648 12189
rect 16590 12121 16602 12155
rect 16636 12121 16648 12155
rect 16590 12087 16648 12121
rect 16590 12053 16602 12087
rect 16636 12053 16648 12087
rect 16590 12019 16648 12053
rect 16590 11985 16602 12019
rect 16636 11985 16648 12019
rect 16590 11951 16648 11985
rect 16590 11917 16602 11951
rect 16636 11917 16648 11951
rect 16590 11883 16648 11917
rect 16590 11849 16602 11883
rect 16636 11849 16648 11883
rect 16590 11815 16648 11849
rect 16590 11781 16602 11815
rect 16636 11781 16648 11815
rect 16590 11747 16648 11781
rect 16590 11713 16602 11747
rect 16636 11713 16648 11747
rect 16590 11679 16648 11713
rect 16590 11645 16602 11679
rect 16636 11645 16648 11679
rect 16590 11611 16648 11645
rect 16590 11577 16602 11611
rect 16636 11577 16648 11611
rect 16590 11543 16648 11577
rect 16590 11509 16602 11543
rect 16636 11509 16648 11543
rect 16590 11475 16648 11509
rect 16590 11441 16602 11475
rect 16636 11441 16648 11475
rect 16590 11407 16648 11441
rect 16590 11373 16602 11407
rect 16636 11373 16648 11407
rect 16590 11339 16648 11373
rect 16590 11305 16602 11339
rect 16636 11305 16648 11339
rect 16590 11271 16648 11305
rect 16590 11237 16602 11271
rect 16636 11237 16648 11271
rect 16590 11203 16648 11237
rect 16590 11169 16602 11203
rect 16636 11169 16648 11203
rect 16590 11135 16648 11169
rect 16590 11101 16602 11135
rect 16636 11101 16648 11135
rect 16590 11070 16648 11101
rect 16678 13039 16736 13070
rect 16678 13005 16690 13039
rect 16724 13005 16736 13039
rect 16678 12971 16736 13005
rect 16678 12937 16690 12971
rect 16724 12937 16736 12971
rect 16678 12903 16736 12937
rect 16678 12869 16690 12903
rect 16724 12869 16736 12903
rect 16678 12835 16736 12869
rect 16678 12801 16690 12835
rect 16724 12801 16736 12835
rect 16678 12767 16736 12801
rect 16678 12733 16690 12767
rect 16724 12733 16736 12767
rect 16678 12699 16736 12733
rect 16678 12665 16690 12699
rect 16724 12665 16736 12699
rect 16678 12631 16736 12665
rect 16678 12597 16690 12631
rect 16724 12597 16736 12631
rect 16678 12563 16736 12597
rect 16678 12529 16690 12563
rect 16724 12529 16736 12563
rect 16678 12495 16736 12529
rect 16678 12461 16690 12495
rect 16724 12461 16736 12495
rect 16678 12427 16736 12461
rect 16678 12393 16690 12427
rect 16724 12393 16736 12427
rect 16678 12359 16736 12393
rect 16678 12325 16690 12359
rect 16724 12325 16736 12359
rect 16678 12291 16736 12325
rect 16678 12257 16690 12291
rect 16724 12257 16736 12291
rect 16678 12223 16736 12257
rect 16678 12189 16690 12223
rect 16724 12189 16736 12223
rect 16678 12155 16736 12189
rect 16678 12121 16690 12155
rect 16724 12121 16736 12155
rect 16678 12087 16736 12121
rect 16678 12053 16690 12087
rect 16724 12053 16736 12087
rect 16678 12019 16736 12053
rect 16678 11985 16690 12019
rect 16724 11985 16736 12019
rect 16678 11951 16736 11985
rect 16678 11917 16690 11951
rect 16724 11917 16736 11951
rect 16678 11883 16736 11917
rect 16678 11849 16690 11883
rect 16724 11849 16736 11883
rect 16678 11815 16736 11849
rect 16678 11781 16690 11815
rect 16724 11781 16736 11815
rect 16678 11747 16736 11781
rect 16678 11713 16690 11747
rect 16724 11713 16736 11747
rect 16678 11679 16736 11713
rect 16678 11645 16690 11679
rect 16724 11645 16736 11679
rect 16678 11611 16736 11645
rect 16678 11577 16690 11611
rect 16724 11577 16736 11611
rect 16678 11543 16736 11577
rect 16678 11509 16690 11543
rect 16724 11509 16736 11543
rect 16678 11475 16736 11509
rect 16678 11441 16690 11475
rect 16724 11441 16736 11475
rect 16678 11407 16736 11441
rect 16678 11373 16690 11407
rect 16724 11373 16736 11407
rect 16678 11339 16736 11373
rect 16678 11305 16690 11339
rect 16724 11305 16736 11339
rect 16678 11271 16736 11305
rect 16678 11237 16690 11271
rect 16724 11237 16736 11271
rect 16678 11203 16736 11237
rect 16678 11169 16690 11203
rect 16724 11169 16736 11203
rect 16678 11135 16736 11169
rect 16678 11101 16690 11135
rect 16724 11101 16736 11135
rect 16678 11070 16736 11101
rect 16766 13039 16824 13070
rect 16766 13005 16778 13039
rect 16812 13005 16824 13039
rect 16766 12971 16824 13005
rect 16766 12937 16778 12971
rect 16812 12937 16824 12971
rect 16766 12903 16824 12937
rect 16766 12869 16778 12903
rect 16812 12869 16824 12903
rect 16766 12835 16824 12869
rect 16766 12801 16778 12835
rect 16812 12801 16824 12835
rect 16766 12767 16824 12801
rect 16766 12733 16778 12767
rect 16812 12733 16824 12767
rect 16766 12699 16824 12733
rect 16766 12665 16778 12699
rect 16812 12665 16824 12699
rect 16766 12631 16824 12665
rect 16766 12597 16778 12631
rect 16812 12597 16824 12631
rect 16766 12563 16824 12597
rect 16766 12529 16778 12563
rect 16812 12529 16824 12563
rect 16766 12495 16824 12529
rect 16766 12461 16778 12495
rect 16812 12461 16824 12495
rect 16766 12427 16824 12461
rect 16766 12393 16778 12427
rect 16812 12393 16824 12427
rect 16766 12359 16824 12393
rect 16766 12325 16778 12359
rect 16812 12325 16824 12359
rect 16766 12291 16824 12325
rect 16766 12257 16778 12291
rect 16812 12257 16824 12291
rect 16766 12223 16824 12257
rect 16766 12189 16778 12223
rect 16812 12189 16824 12223
rect 16766 12155 16824 12189
rect 16766 12121 16778 12155
rect 16812 12121 16824 12155
rect 16766 12087 16824 12121
rect 16766 12053 16778 12087
rect 16812 12053 16824 12087
rect 16766 12019 16824 12053
rect 16766 11985 16778 12019
rect 16812 11985 16824 12019
rect 16766 11951 16824 11985
rect 16766 11917 16778 11951
rect 16812 11917 16824 11951
rect 16766 11883 16824 11917
rect 16766 11849 16778 11883
rect 16812 11849 16824 11883
rect 16766 11815 16824 11849
rect 16766 11781 16778 11815
rect 16812 11781 16824 11815
rect 16766 11747 16824 11781
rect 16766 11713 16778 11747
rect 16812 11713 16824 11747
rect 16766 11679 16824 11713
rect 16766 11645 16778 11679
rect 16812 11645 16824 11679
rect 16766 11611 16824 11645
rect 16766 11577 16778 11611
rect 16812 11577 16824 11611
rect 16766 11543 16824 11577
rect 16766 11509 16778 11543
rect 16812 11509 16824 11543
rect 16766 11475 16824 11509
rect 16766 11441 16778 11475
rect 16812 11441 16824 11475
rect 16766 11407 16824 11441
rect 16766 11373 16778 11407
rect 16812 11373 16824 11407
rect 16766 11339 16824 11373
rect 16766 11305 16778 11339
rect 16812 11305 16824 11339
rect 16766 11271 16824 11305
rect 16766 11237 16778 11271
rect 16812 11237 16824 11271
rect 16766 11203 16824 11237
rect 16766 11169 16778 11203
rect 16812 11169 16824 11203
rect 16766 11135 16824 11169
rect 16766 11101 16778 11135
rect 16812 11101 16824 11135
rect 16766 11070 16824 11101
rect 16854 13039 16912 13070
rect 16854 13005 16866 13039
rect 16900 13005 16912 13039
rect 16854 12971 16912 13005
rect 16854 12937 16866 12971
rect 16900 12937 16912 12971
rect 16854 12903 16912 12937
rect 16854 12869 16866 12903
rect 16900 12869 16912 12903
rect 16854 12835 16912 12869
rect 16854 12801 16866 12835
rect 16900 12801 16912 12835
rect 16854 12767 16912 12801
rect 16854 12733 16866 12767
rect 16900 12733 16912 12767
rect 16854 12699 16912 12733
rect 16854 12665 16866 12699
rect 16900 12665 16912 12699
rect 16854 12631 16912 12665
rect 16854 12597 16866 12631
rect 16900 12597 16912 12631
rect 16854 12563 16912 12597
rect 16854 12529 16866 12563
rect 16900 12529 16912 12563
rect 16854 12495 16912 12529
rect 16854 12461 16866 12495
rect 16900 12461 16912 12495
rect 16854 12427 16912 12461
rect 16854 12393 16866 12427
rect 16900 12393 16912 12427
rect 16854 12359 16912 12393
rect 16854 12325 16866 12359
rect 16900 12325 16912 12359
rect 16854 12291 16912 12325
rect 16854 12257 16866 12291
rect 16900 12257 16912 12291
rect 16854 12223 16912 12257
rect 16854 12189 16866 12223
rect 16900 12189 16912 12223
rect 16854 12155 16912 12189
rect 16854 12121 16866 12155
rect 16900 12121 16912 12155
rect 16854 12087 16912 12121
rect 16854 12053 16866 12087
rect 16900 12053 16912 12087
rect 16854 12019 16912 12053
rect 16854 11985 16866 12019
rect 16900 11985 16912 12019
rect 16854 11951 16912 11985
rect 16854 11917 16866 11951
rect 16900 11917 16912 11951
rect 16854 11883 16912 11917
rect 16854 11849 16866 11883
rect 16900 11849 16912 11883
rect 16854 11815 16912 11849
rect 16854 11781 16866 11815
rect 16900 11781 16912 11815
rect 16854 11747 16912 11781
rect 16854 11713 16866 11747
rect 16900 11713 16912 11747
rect 16854 11679 16912 11713
rect 16854 11645 16866 11679
rect 16900 11645 16912 11679
rect 16854 11611 16912 11645
rect 16854 11577 16866 11611
rect 16900 11577 16912 11611
rect 16854 11543 16912 11577
rect 16854 11509 16866 11543
rect 16900 11509 16912 11543
rect 16854 11475 16912 11509
rect 16854 11441 16866 11475
rect 16900 11441 16912 11475
rect 16854 11407 16912 11441
rect 16854 11373 16866 11407
rect 16900 11373 16912 11407
rect 16854 11339 16912 11373
rect 16854 11305 16866 11339
rect 16900 11305 16912 11339
rect 16854 11271 16912 11305
rect 16854 11237 16866 11271
rect 16900 11237 16912 11271
rect 16854 11203 16912 11237
rect 16854 11169 16866 11203
rect 16900 11169 16912 11203
rect 16854 11135 16912 11169
rect 16854 11101 16866 11135
rect 16900 11101 16912 11135
rect 16854 11070 16912 11101
rect 16942 13039 17000 13070
rect 16942 13005 16954 13039
rect 16988 13005 17000 13039
rect 16942 12971 17000 13005
rect 16942 12937 16954 12971
rect 16988 12937 17000 12971
rect 16942 12903 17000 12937
rect 16942 12869 16954 12903
rect 16988 12869 17000 12903
rect 16942 12835 17000 12869
rect 16942 12801 16954 12835
rect 16988 12801 17000 12835
rect 16942 12767 17000 12801
rect 16942 12733 16954 12767
rect 16988 12733 17000 12767
rect 16942 12699 17000 12733
rect 16942 12665 16954 12699
rect 16988 12665 17000 12699
rect 16942 12631 17000 12665
rect 16942 12597 16954 12631
rect 16988 12597 17000 12631
rect 16942 12563 17000 12597
rect 16942 12529 16954 12563
rect 16988 12529 17000 12563
rect 16942 12495 17000 12529
rect 16942 12461 16954 12495
rect 16988 12461 17000 12495
rect 16942 12427 17000 12461
rect 16942 12393 16954 12427
rect 16988 12393 17000 12427
rect 16942 12359 17000 12393
rect 16942 12325 16954 12359
rect 16988 12325 17000 12359
rect 16942 12291 17000 12325
rect 16942 12257 16954 12291
rect 16988 12257 17000 12291
rect 16942 12223 17000 12257
rect 16942 12189 16954 12223
rect 16988 12189 17000 12223
rect 16942 12155 17000 12189
rect 16942 12121 16954 12155
rect 16988 12121 17000 12155
rect 16942 12087 17000 12121
rect 16942 12053 16954 12087
rect 16988 12053 17000 12087
rect 16942 12019 17000 12053
rect 16942 11985 16954 12019
rect 16988 11985 17000 12019
rect 16942 11951 17000 11985
rect 16942 11917 16954 11951
rect 16988 11917 17000 11951
rect 16942 11883 17000 11917
rect 16942 11849 16954 11883
rect 16988 11849 17000 11883
rect 16942 11815 17000 11849
rect 16942 11781 16954 11815
rect 16988 11781 17000 11815
rect 16942 11747 17000 11781
rect 16942 11713 16954 11747
rect 16988 11713 17000 11747
rect 16942 11679 17000 11713
rect 16942 11645 16954 11679
rect 16988 11645 17000 11679
rect 16942 11611 17000 11645
rect 16942 11577 16954 11611
rect 16988 11577 17000 11611
rect 16942 11543 17000 11577
rect 16942 11509 16954 11543
rect 16988 11509 17000 11543
rect 16942 11475 17000 11509
rect 16942 11441 16954 11475
rect 16988 11441 17000 11475
rect 16942 11407 17000 11441
rect 16942 11373 16954 11407
rect 16988 11373 17000 11407
rect 16942 11339 17000 11373
rect 16942 11305 16954 11339
rect 16988 11305 17000 11339
rect 16942 11271 17000 11305
rect 16942 11237 16954 11271
rect 16988 11237 17000 11271
rect 16942 11203 17000 11237
rect 16942 11169 16954 11203
rect 16988 11169 17000 11203
rect 16942 11135 17000 11169
rect 16942 11101 16954 11135
rect 16988 11101 17000 11135
rect 16942 11070 17000 11101
rect 17030 13039 17088 13070
rect 17030 13005 17042 13039
rect 17076 13005 17088 13039
rect 17030 12971 17088 13005
rect 17030 12937 17042 12971
rect 17076 12937 17088 12971
rect 17030 12903 17088 12937
rect 17030 12869 17042 12903
rect 17076 12869 17088 12903
rect 17030 12835 17088 12869
rect 17030 12801 17042 12835
rect 17076 12801 17088 12835
rect 17030 12767 17088 12801
rect 17030 12733 17042 12767
rect 17076 12733 17088 12767
rect 17030 12699 17088 12733
rect 17030 12665 17042 12699
rect 17076 12665 17088 12699
rect 17030 12631 17088 12665
rect 17030 12597 17042 12631
rect 17076 12597 17088 12631
rect 17030 12563 17088 12597
rect 17030 12529 17042 12563
rect 17076 12529 17088 12563
rect 17030 12495 17088 12529
rect 17030 12461 17042 12495
rect 17076 12461 17088 12495
rect 17030 12427 17088 12461
rect 17030 12393 17042 12427
rect 17076 12393 17088 12427
rect 17030 12359 17088 12393
rect 17030 12325 17042 12359
rect 17076 12325 17088 12359
rect 17030 12291 17088 12325
rect 17030 12257 17042 12291
rect 17076 12257 17088 12291
rect 17030 12223 17088 12257
rect 17030 12189 17042 12223
rect 17076 12189 17088 12223
rect 17030 12155 17088 12189
rect 17030 12121 17042 12155
rect 17076 12121 17088 12155
rect 17030 12087 17088 12121
rect 17030 12053 17042 12087
rect 17076 12053 17088 12087
rect 17030 12019 17088 12053
rect 17030 11985 17042 12019
rect 17076 11985 17088 12019
rect 17030 11951 17088 11985
rect 17030 11917 17042 11951
rect 17076 11917 17088 11951
rect 17030 11883 17088 11917
rect 17030 11849 17042 11883
rect 17076 11849 17088 11883
rect 17030 11815 17088 11849
rect 17030 11781 17042 11815
rect 17076 11781 17088 11815
rect 17030 11747 17088 11781
rect 17030 11713 17042 11747
rect 17076 11713 17088 11747
rect 17030 11679 17088 11713
rect 17030 11645 17042 11679
rect 17076 11645 17088 11679
rect 17030 11611 17088 11645
rect 17030 11577 17042 11611
rect 17076 11577 17088 11611
rect 17030 11543 17088 11577
rect 17030 11509 17042 11543
rect 17076 11509 17088 11543
rect 17030 11475 17088 11509
rect 17030 11441 17042 11475
rect 17076 11441 17088 11475
rect 17030 11407 17088 11441
rect 17030 11373 17042 11407
rect 17076 11373 17088 11407
rect 17030 11339 17088 11373
rect 17030 11305 17042 11339
rect 17076 11305 17088 11339
rect 17030 11271 17088 11305
rect 17030 11237 17042 11271
rect 17076 11237 17088 11271
rect 17030 11203 17088 11237
rect 17030 11169 17042 11203
rect 17076 11169 17088 11203
rect 17030 11135 17088 11169
rect 17030 11101 17042 11135
rect 17076 11101 17088 11135
rect 17030 11070 17088 11101
rect 17118 13039 17176 13070
rect 17118 13005 17130 13039
rect 17164 13005 17176 13039
rect 17118 12971 17176 13005
rect 17118 12937 17130 12971
rect 17164 12937 17176 12971
rect 17118 12903 17176 12937
rect 17118 12869 17130 12903
rect 17164 12869 17176 12903
rect 17118 12835 17176 12869
rect 17118 12801 17130 12835
rect 17164 12801 17176 12835
rect 17118 12767 17176 12801
rect 17118 12733 17130 12767
rect 17164 12733 17176 12767
rect 17118 12699 17176 12733
rect 17118 12665 17130 12699
rect 17164 12665 17176 12699
rect 17118 12631 17176 12665
rect 17118 12597 17130 12631
rect 17164 12597 17176 12631
rect 17118 12563 17176 12597
rect 17118 12529 17130 12563
rect 17164 12529 17176 12563
rect 17118 12495 17176 12529
rect 17118 12461 17130 12495
rect 17164 12461 17176 12495
rect 17118 12427 17176 12461
rect 17118 12393 17130 12427
rect 17164 12393 17176 12427
rect 17118 12359 17176 12393
rect 17118 12325 17130 12359
rect 17164 12325 17176 12359
rect 17118 12291 17176 12325
rect 17118 12257 17130 12291
rect 17164 12257 17176 12291
rect 17118 12223 17176 12257
rect 17118 12189 17130 12223
rect 17164 12189 17176 12223
rect 17118 12155 17176 12189
rect 17118 12121 17130 12155
rect 17164 12121 17176 12155
rect 17118 12087 17176 12121
rect 17118 12053 17130 12087
rect 17164 12053 17176 12087
rect 17118 12019 17176 12053
rect 17118 11985 17130 12019
rect 17164 11985 17176 12019
rect 17118 11951 17176 11985
rect 17118 11917 17130 11951
rect 17164 11917 17176 11951
rect 17118 11883 17176 11917
rect 17118 11849 17130 11883
rect 17164 11849 17176 11883
rect 17118 11815 17176 11849
rect 17118 11781 17130 11815
rect 17164 11781 17176 11815
rect 17118 11747 17176 11781
rect 17118 11713 17130 11747
rect 17164 11713 17176 11747
rect 17118 11679 17176 11713
rect 17118 11645 17130 11679
rect 17164 11645 17176 11679
rect 17118 11611 17176 11645
rect 17118 11577 17130 11611
rect 17164 11577 17176 11611
rect 17118 11543 17176 11577
rect 17118 11509 17130 11543
rect 17164 11509 17176 11543
rect 17118 11475 17176 11509
rect 17118 11441 17130 11475
rect 17164 11441 17176 11475
rect 17118 11407 17176 11441
rect 17118 11373 17130 11407
rect 17164 11373 17176 11407
rect 17118 11339 17176 11373
rect 17118 11305 17130 11339
rect 17164 11305 17176 11339
rect 17118 11271 17176 11305
rect 17118 11237 17130 11271
rect 17164 11237 17176 11271
rect 17118 11203 17176 11237
rect 17118 11169 17130 11203
rect 17164 11169 17176 11203
rect 17118 11135 17176 11169
rect 17118 11101 17130 11135
rect 17164 11101 17176 11135
rect 17118 11070 17176 11101
rect 17206 13039 17264 13070
rect 17206 13005 17218 13039
rect 17252 13005 17264 13039
rect 17206 12971 17264 13005
rect 17206 12937 17218 12971
rect 17252 12937 17264 12971
rect 17206 12903 17264 12937
rect 17206 12869 17218 12903
rect 17252 12869 17264 12903
rect 17206 12835 17264 12869
rect 17206 12801 17218 12835
rect 17252 12801 17264 12835
rect 17206 12767 17264 12801
rect 17206 12733 17218 12767
rect 17252 12733 17264 12767
rect 17206 12699 17264 12733
rect 17206 12665 17218 12699
rect 17252 12665 17264 12699
rect 17206 12631 17264 12665
rect 17206 12597 17218 12631
rect 17252 12597 17264 12631
rect 17206 12563 17264 12597
rect 17206 12529 17218 12563
rect 17252 12529 17264 12563
rect 17206 12495 17264 12529
rect 17206 12461 17218 12495
rect 17252 12461 17264 12495
rect 17206 12427 17264 12461
rect 17206 12393 17218 12427
rect 17252 12393 17264 12427
rect 17206 12359 17264 12393
rect 17206 12325 17218 12359
rect 17252 12325 17264 12359
rect 17206 12291 17264 12325
rect 17206 12257 17218 12291
rect 17252 12257 17264 12291
rect 17206 12223 17264 12257
rect 17206 12189 17218 12223
rect 17252 12189 17264 12223
rect 17206 12155 17264 12189
rect 17206 12121 17218 12155
rect 17252 12121 17264 12155
rect 17206 12087 17264 12121
rect 17206 12053 17218 12087
rect 17252 12053 17264 12087
rect 17206 12019 17264 12053
rect 17206 11985 17218 12019
rect 17252 11985 17264 12019
rect 17206 11951 17264 11985
rect 17206 11917 17218 11951
rect 17252 11917 17264 11951
rect 17206 11883 17264 11917
rect 17206 11849 17218 11883
rect 17252 11849 17264 11883
rect 17206 11815 17264 11849
rect 17206 11781 17218 11815
rect 17252 11781 17264 11815
rect 17206 11747 17264 11781
rect 17206 11713 17218 11747
rect 17252 11713 17264 11747
rect 17206 11679 17264 11713
rect 17206 11645 17218 11679
rect 17252 11645 17264 11679
rect 17206 11611 17264 11645
rect 17206 11577 17218 11611
rect 17252 11577 17264 11611
rect 17206 11543 17264 11577
rect 17206 11509 17218 11543
rect 17252 11509 17264 11543
rect 17206 11475 17264 11509
rect 17206 11441 17218 11475
rect 17252 11441 17264 11475
rect 17206 11407 17264 11441
rect 17206 11373 17218 11407
rect 17252 11373 17264 11407
rect 17206 11339 17264 11373
rect 17206 11305 17218 11339
rect 17252 11305 17264 11339
rect 17206 11271 17264 11305
rect 17206 11237 17218 11271
rect 17252 11237 17264 11271
rect 17206 11203 17264 11237
rect 17206 11169 17218 11203
rect 17252 11169 17264 11203
rect 17206 11135 17264 11169
rect 17206 11101 17218 11135
rect 17252 11101 17264 11135
rect 17206 11070 17264 11101
rect 17294 13039 17352 13070
rect 17294 13005 17306 13039
rect 17340 13005 17352 13039
rect 17294 12971 17352 13005
rect 17294 12937 17306 12971
rect 17340 12937 17352 12971
rect 17294 12903 17352 12937
rect 17294 12869 17306 12903
rect 17340 12869 17352 12903
rect 17294 12835 17352 12869
rect 17294 12801 17306 12835
rect 17340 12801 17352 12835
rect 17294 12767 17352 12801
rect 17294 12733 17306 12767
rect 17340 12733 17352 12767
rect 17294 12699 17352 12733
rect 17294 12665 17306 12699
rect 17340 12665 17352 12699
rect 17294 12631 17352 12665
rect 17294 12597 17306 12631
rect 17340 12597 17352 12631
rect 17294 12563 17352 12597
rect 17294 12529 17306 12563
rect 17340 12529 17352 12563
rect 17294 12495 17352 12529
rect 17294 12461 17306 12495
rect 17340 12461 17352 12495
rect 17294 12427 17352 12461
rect 17294 12393 17306 12427
rect 17340 12393 17352 12427
rect 17294 12359 17352 12393
rect 17294 12325 17306 12359
rect 17340 12325 17352 12359
rect 17294 12291 17352 12325
rect 17294 12257 17306 12291
rect 17340 12257 17352 12291
rect 17294 12223 17352 12257
rect 17294 12189 17306 12223
rect 17340 12189 17352 12223
rect 17294 12155 17352 12189
rect 17294 12121 17306 12155
rect 17340 12121 17352 12155
rect 17294 12087 17352 12121
rect 17294 12053 17306 12087
rect 17340 12053 17352 12087
rect 17294 12019 17352 12053
rect 17294 11985 17306 12019
rect 17340 11985 17352 12019
rect 17294 11951 17352 11985
rect 17294 11917 17306 11951
rect 17340 11917 17352 11951
rect 17294 11883 17352 11917
rect 17294 11849 17306 11883
rect 17340 11849 17352 11883
rect 17294 11815 17352 11849
rect 17294 11781 17306 11815
rect 17340 11781 17352 11815
rect 17294 11747 17352 11781
rect 17294 11713 17306 11747
rect 17340 11713 17352 11747
rect 17294 11679 17352 11713
rect 17294 11645 17306 11679
rect 17340 11645 17352 11679
rect 17294 11611 17352 11645
rect 17294 11577 17306 11611
rect 17340 11577 17352 11611
rect 17294 11543 17352 11577
rect 17294 11509 17306 11543
rect 17340 11509 17352 11543
rect 17294 11475 17352 11509
rect 17294 11441 17306 11475
rect 17340 11441 17352 11475
rect 17294 11407 17352 11441
rect 17294 11373 17306 11407
rect 17340 11373 17352 11407
rect 17294 11339 17352 11373
rect 17294 11305 17306 11339
rect 17340 11305 17352 11339
rect 17294 11271 17352 11305
rect 17294 11237 17306 11271
rect 17340 11237 17352 11271
rect 17294 11203 17352 11237
rect 17294 11169 17306 11203
rect 17340 11169 17352 11203
rect 17294 11135 17352 11169
rect 17294 11101 17306 11135
rect 17340 11101 17352 11135
rect 17294 11070 17352 11101
rect 17382 13039 17440 13070
rect 17382 13005 17394 13039
rect 17428 13005 17440 13039
rect 17382 12971 17440 13005
rect 17382 12937 17394 12971
rect 17428 12937 17440 12971
rect 17382 12903 17440 12937
rect 17382 12869 17394 12903
rect 17428 12869 17440 12903
rect 17382 12835 17440 12869
rect 17382 12801 17394 12835
rect 17428 12801 17440 12835
rect 17382 12767 17440 12801
rect 17382 12733 17394 12767
rect 17428 12733 17440 12767
rect 17382 12699 17440 12733
rect 17382 12665 17394 12699
rect 17428 12665 17440 12699
rect 17382 12631 17440 12665
rect 17382 12597 17394 12631
rect 17428 12597 17440 12631
rect 17382 12563 17440 12597
rect 17382 12529 17394 12563
rect 17428 12529 17440 12563
rect 17382 12495 17440 12529
rect 17382 12461 17394 12495
rect 17428 12461 17440 12495
rect 17382 12427 17440 12461
rect 17382 12393 17394 12427
rect 17428 12393 17440 12427
rect 17382 12359 17440 12393
rect 17382 12325 17394 12359
rect 17428 12325 17440 12359
rect 17382 12291 17440 12325
rect 17382 12257 17394 12291
rect 17428 12257 17440 12291
rect 17382 12223 17440 12257
rect 17382 12189 17394 12223
rect 17428 12189 17440 12223
rect 17382 12155 17440 12189
rect 17382 12121 17394 12155
rect 17428 12121 17440 12155
rect 17382 12087 17440 12121
rect 17382 12053 17394 12087
rect 17428 12053 17440 12087
rect 17382 12019 17440 12053
rect 17382 11985 17394 12019
rect 17428 11985 17440 12019
rect 17382 11951 17440 11985
rect 17382 11917 17394 11951
rect 17428 11917 17440 11951
rect 17382 11883 17440 11917
rect 17382 11849 17394 11883
rect 17428 11849 17440 11883
rect 17382 11815 17440 11849
rect 17382 11781 17394 11815
rect 17428 11781 17440 11815
rect 17382 11747 17440 11781
rect 17382 11713 17394 11747
rect 17428 11713 17440 11747
rect 17382 11679 17440 11713
rect 17382 11645 17394 11679
rect 17428 11645 17440 11679
rect 17382 11611 17440 11645
rect 17382 11577 17394 11611
rect 17428 11577 17440 11611
rect 17382 11543 17440 11577
rect 17382 11509 17394 11543
rect 17428 11509 17440 11543
rect 17382 11475 17440 11509
rect 17382 11441 17394 11475
rect 17428 11441 17440 11475
rect 17382 11407 17440 11441
rect 17382 11373 17394 11407
rect 17428 11373 17440 11407
rect 17382 11339 17440 11373
rect 17382 11305 17394 11339
rect 17428 11305 17440 11339
rect 17382 11271 17440 11305
rect 17382 11237 17394 11271
rect 17428 11237 17440 11271
rect 17382 11203 17440 11237
rect 17382 11169 17394 11203
rect 17428 11169 17440 11203
rect 17382 11135 17440 11169
rect 17382 11101 17394 11135
rect 17428 11101 17440 11135
rect 17382 11070 17440 11101
rect 17470 13039 17528 13070
rect 17470 13005 17482 13039
rect 17516 13005 17528 13039
rect 17470 12971 17528 13005
rect 17470 12937 17482 12971
rect 17516 12937 17528 12971
rect 17470 12903 17528 12937
rect 17470 12869 17482 12903
rect 17516 12869 17528 12903
rect 17470 12835 17528 12869
rect 17470 12801 17482 12835
rect 17516 12801 17528 12835
rect 17470 12767 17528 12801
rect 17470 12733 17482 12767
rect 17516 12733 17528 12767
rect 17470 12699 17528 12733
rect 17470 12665 17482 12699
rect 17516 12665 17528 12699
rect 17470 12631 17528 12665
rect 17470 12597 17482 12631
rect 17516 12597 17528 12631
rect 17470 12563 17528 12597
rect 17470 12529 17482 12563
rect 17516 12529 17528 12563
rect 17470 12495 17528 12529
rect 17470 12461 17482 12495
rect 17516 12461 17528 12495
rect 17470 12427 17528 12461
rect 17470 12393 17482 12427
rect 17516 12393 17528 12427
rect 17470 12359 17528 12393
rect 17470 12325 17482 12359
rect 17516 12325 17528 12359
rect 17470 12291 17528 12325
rect 17470 12257 17482 12291
rect 17516 12257 17528 12291
rect 17470 12223 17528 12257
rect 17470 12189 17482 12223
rect 17516 12189 17528 12223
rect 17470 12155 17528 12189
rect 17470 12121 17482 12155
rect 17516 12121 17528 12155
rect 17470 12087 17528 12121
rect 17470 12053 17482 12087
rect 17516 12053 17528 12087
rect 17470 12019 17528 12053
rect 17470 11985 17482 12019
rect 17516 11985 17528 12019
rect 17470 11951 17528 11985
rect 17470 11917 17482 11951
rect 17516 11917 17528 11951
rect 17470 11883 17528 11917
rect 17470 11849 17482 11883
rect 17516 11849 17528 11883
rect 17470 11815 17528 11849
rect 17470 11781 17482 11815
rect 17516 11781 17528 11815
rect 17470 11747 17528 11781
rect 17470 11713 17482 11747
rect 17516 11713 17528 11747
rect 17470 11679 17528 11713
rect 17470 11645 17482 11679
rect 17516 11645 17528 11679
rect 17470 11611 17528 11645
rect 17470 11577 17482 11611
rect 17516 11577 17528 11611
rect 17470 11543 17528 11577
rect 17470 11509 17482 11543
rect 17516 11509 17528 11543
rect 17470 11475 17528 11509
rect 17470 11441 17482 11475
rect 17516 11441 17528 11475
rect 17470 11407 17528 11441
rect 17470 11373 17482 11407
rect 17516 11373 17528 11407
rect 17470 11339 17528 11373
rect 17470 11305 17482 11339
rect 17516 11305 17528 11339
rect 17470 11271 17528 11305
rect 17470 11237 17482 11271
rect 17516 11237 17528 11271
rect 17470 11203 17528 11237
rect 17470 11169 17482 11203
rect 17516 11169 17528 11203
rect 17470 11135 17528 11169
rect 17470 11101 17482 11135
rect 17516 11101 17528 11135
rect 17470 11070 17528 11101
<< pdiff >>
rect 15818 23158 15880 23189
rect 15818 23124 15830 23158
rect 15864 23124 15880 23158
rect 15818 23090 15880 23124
rect 15818 23056 15830 23090
rect 15864 23056 15880 23090
rect 15818 23022 15880 23056
rect 15818 22988 15830 23022
rect 15864 22988 15880 23022
rect 15818 22954 15880 22988
rect 15818 22920 15830 22954
rect 15864 22920 15880 22954
rect 15818 22886 15880 22920
rect 15818 22852 15830 22886
rect 15864 22852 15880 22886
rect 15818 22818 15880 22852
rect 15818 22784 15830 22818
rect 15864 22784 15880 22818
rect 15818 22750 15880 22784
rect 15818 22716 15830 22750
rect 15864 22716 15880 22750
rect 15818 22682 15880 22716
rect 15818 22648 15830 22682
rect 15864 22648 15880 22682
rect 15818 22614 15880 22648
rect 15818 22580 15830 22614
rect 15864 22580 15880 22614
rect 15818 22546 15880 22580
rect 15818 22512 15830 22546
rect 15864 22512 15880 22546
rect 15818 22478 15880 22512
rect 15818 22444 15830 22478
rect 15864 22444 15880 22478
rect 15818 22410 15880 22444
rect 15818 22376 15830 22410
rect 15864 22376 15880 22410
rect 15818 22342 15880 22376
rect 15818 22308 15830 22342
rect 15864 22308 15880 22342
rect 15818 22274 15880 22308
rect 15818 22240 15830 22274
rect 15864 22240 15880 22274
rect 15818 22206 15880 22240
rect 15818 22172 15830 22206
rect 15864 22172 15880 22206
rect 15818 22138 15880 22172
rect 15818 22104 15830 22138
rect 15864 22104 15880 22138
rect 15818 22070 15880 22104
rect 15818 22036 15830 22070
rect 15864 22036 15880 22070
rect 15818 22002 15880 22036
rect 15818 21968 15830 22002
rect 15864 21968 15880 22002
rect 15818 21934 15880 21968
rect 15818 21900 15830 21934
rect 15864 21900 15880 21934
rect 15818 21866 15880 21900
rect 15818 21832 15830 21866
rect 15864 21832 15880 21866
rect 15818 21798 15880 21832
rect 15818 21764 15830 21798
rect 15864 21764 15880 21798
rect 15818 21730 15880 21764
rect 15818 21696 15830 21730
rect 15864 21696 15880 21730
rect 15818 21662 15880 21696
rect 15818 21628 15830 21662
rect 15864 21628 15880 21662
rect 15818 21594 15880 21628
rect 15818 21560 15830 21594
rect 15864 21560 15880 21594
rect 15818 21526 15880 21560
rect 15818 21492 15830 21526
rect 15864 21492 15880 21526
rect 15818 21458 15880 21492
rect 15818 21424 15830 21458
rect 15864 21424 15880 21458
rect 15818 21390 15880 21424
rect 15818 21356 15830 21390
rect 15864 21356 15880 21390
rect 15818 21322 15880 21356
rect 15818 21288 15830 21322
rect 15864 21288 15880 21322
rect 15818 21254 15880 21288
rect 15818 21220 15830 21254
rect 15864 21220 15880 21254
rect 15818 21189 15880 21220
rect 15910 23158 15976 23189
rect 15910 23124 15926 23158
rect 15960 23124 15976 23158
rect 15910 23090 15976 23124
rect 15910 23056 15926 23090
rect 15960 23056 15976 23090
rect 15910 23022 15976 23056
rect 15910 22988 15926 23022
rect 15960 22988 15976 23022
rect 15910 22954 15976 22988
rect 15910 22920 15926 22954
rect 15960 22920 15976 22954
rect 15910 22886 15976 22920
rect 15910 22852 15926 22886
rect 15960 22852 15976 22886
rect 15910 22818 15976 22852
rect 15910 22784 15926 22818
rect 15960 22784 15976 22818
rect 15910 22750 15976 22784
rect 15910 22716 15926 22750
rect 15960 22716 15976 22750
rect 15910 22682 15976 22716
rect 15910 22648 15926 22682
rect 15960 22648 15976 22682
rect 15910 22614 15976 22648
rect 15910 22580 15926 22614
rect 15960 22580 15976 22614
rect 15910 22546 15976 22580
rect 15910 22512 15926 22546
rect 15960 22512 15976 22546
rect 15910 22478 15976 22512
rect 15910 22444 15926 22478
rect 15960 22444 15976 22478
rect 15910 22410 15976 22444
rect 15910 22376 15926 22410
rect 15960 22376 15976 22410
rect 15910 22342 15976 22376
rect 15910 22308 15926 22342
rect 15960 22308 15976 22342
rect 15910 22274 15976 22308
rect 15910 22240 15926 22274
rect 15960 22240 15976 22274
rect 15910 22206 15976 22240
rect 15910 22172 15926 22206
rect 15960 22172 15976 22206
rect 15910 22138 15976 22172
rect 15910 22104 15926 22138
rect 15960 22104 15976 22138
rect 15910 22070 15976 22104
rect 15910 22036 15926 22070
rect 15960 22036 15976 22070
rect 15910 22002 15976 22036
rect 15910 21968 15926 22002
rect 15960 21968 15976 22002
rect 15910 21934 15976 21968
rect 15910 21900 15926 21934
rect 15960 21900 15976 21934
rect 15910 21866 15976 21900
rect 15910 21832 15926 21866
rect 15960 21832 15976 21866
rect 15910 21798 15976 21832
rect 15910 21764 15926 21798
rect 15960 21764 15976 21798
rect 15910 21730 15976 21764
rect 15910 21696 15926 21730
rect 15960 21696 15976 21730
rect 15910 21662 15976 21696
rect 15910 21628 15926 21662
rect 15960 21628 15976 21662
rect 15910 21594 15976 21628
rect 15910 21560 15926 21594
rect 15960 21560 15976 21594
rect 15910 21526 15976 21560
rect 15910 21492 15926 21526
rect 15960 21492 15976 21526
rect 15910 21458 15976 21492
rect 15910 21424 15926 21458
rect 15960 21424 15976 21458
rect 15910 21390 15976 21424
rect 15910 21356 15926 21390
rect 15960 21356 15976 21390
rect 15910 21322 15976 21356
rect 15910 21288 15926 21322
rect 15960 21288 15976 21322
rect 15910 21254 15976 21288
rect 15910 21220 15926 21254
rect 15960 21220 15976 21254
rect 15910 21189 15976 21220
rect 16006 23158 16072 23189
rect 16006 23124 16022 23158
rect 16056 23124 16072 23158
rect 16006 23090 16072 23124
rect 16006 23056 16022 23090
rect 16056 23056 16072 23090
rect 16006 23022 16072 23056
rect 16006 22988 16022 23022
rect 16056 22988 16072 23022
rect 16006 22954 16072 22988
rect 16006 22920 16022 22954
rect 16056 22920 16072 22954
rect 16006 22886 16072 22920
rect 16006 22852 16022 22886
rect 16056 22852 16072 22886
rect 16006 22818 16072 22852
rect 16006 22784 16022 22818
rect 16056 22784 16072 22818
rect 16006 22750 16072 22784
rect 16006 22716 16022 22750
rect 16056 22716 16072 22750
rect 16006 22682 16072 22716
rect 16006 22648 16022 22682
rect 16056 22648 16072 22682
rect 16006 22614 16072 22648
rect 16006 22580 16022 22614
rect 16056 22580 16072 22614
rect 16006 22546 16072 22580
rect 16006 22512 16022 22546
rect 16056 22512 16072 22546
rect 16006 22478 16072 22512
rect 16006 22444 16022 22478
rect 16056 22444 16072 22478
rect 16006 22410 16072 22444
rect 16006 22376 16022 22410
rect 16056 22376 16072 22410
rect 16006 22342 16072 22376
rect 16006 22308 16022 22342
rect 16056 22308 16072 22342
rect 16006 22274 16072 22308
rect 16006 22240 16022 22274
rect 16056 22240 16072 22274
rect 16006 22206 16072 22240
rect 16006 22172 16022 22206
rect 16056 22172 16072 22206
rect 16006 22138 16072 22172
rect 16006 22104 16022 22138
rect 16056 22104 16072 22138
rect 16006 22070 16072 22104
rect 16006 22036 16022 22070
rect 16056 22036 16072 22070
rect 16006 22002 16072 22036
rect 16006 21968 16022 22002
rect 16056 21968 16072 22002
rect 16006 21934 16072 21968
rect 16006 21900 16022 21934
rect 16056 21900 16072 21934
rect 16006 21866 16072 21900
rect 16006 21832 16022 21866
rect 16056 21832 16072 21866
rect 16006 21798 16072 21832
rect 16006 21764 16022 21798
rect 16056 21764 16072 21798
rect 16006 21730 16072 21764
rect 16006 21696 16022 21730
rect 16056 21696 16072 21730
rect 16006 21662 16072 21696
rect 16006 21628 16022 21662
rect 16056 21628 16072 21662
rect 16006 21594 16072 21628
rect 16006 21560 16022 21594
rect 16056 21560 16072 21594
rect 16006 21526 16072 21560
rect 16006 21492 16022 21526
rect 16056 21492 16072 21526
rect 16006 21458 16072 21492
rect 16006 21424 16022 21458
rect 16056 21424 16072 21458
rect 16006 21390 16072 21424
rect 16006 21356 16022 21390
rect 16056 21356 16072 21390
rect 16006 21322 16072 21356
rect 16006 21288 16022 21322
rect 16056 21288 16072 21322
rect 16006 21254 16072 21288
rect 16006 21220 16022 21254
rect 16056 21220 16072 21254
rect 16006 21189 16072 21220
rect 16102 23158 16164 23189
rect 16102 23124 16118 23158
rect 16152 23124 16164 23158
rect 16102 23090 16164 23124
rect 16102 23056 16118 23090
rect 16152 23056 16164 23090
rect 16102 23022 16164 23056
rect 16102 22988 16118 23022
rect 16152 22988 16164 23022
rect 16102 22954 16164 22988
rect 16102 22920 16118 22954
rect 16152 22920 16164 22954
rect 16102 22886 16164 22920
rect 16102 22852 16118 22886
rect 16152 22852 16164 22886
rect 16102 22818 16164 22852
rect 16102 22784 16118 22818
rect 16152 22784 16164 22818
rect 16102 22750 16164 22784
rect 16102 22716 16118 22750
rect 16152 22716 16164 22750
rect 16102 22682 16164 22716
rect 16102 22648 16118 22682
rect 16152 22648 16164 22682
rect 16102 22614 16164 22648
rect 16102 22580 16118 22614
rect 16152 22580 16164 22614
rect 16102 22546 16164 22580
rect 16102 22512 16118 22546
rect 16152 22512 16164 22546
rect 16102 22478 16164 22512
rect 16102 22444 16118 22478
rect 16152 22444 16164 22478
rect 16102 22410 16164 22444
rect 16102 22376 16118 22410
rect 16152 22376 16164 22410
rect 16102 22342 16164 22376
rect 16102 22308 16118 22342
rect 16152 22308 16164 22342
rect 16102 22274 16164 22308
rect 16102 22240 16118 22274
rect 16152 22240 16164 22274
rect 16102 22206 16164 22240
rect 16102 22172 16118 22206
rect 16152 22172 16164 22206
rect 16102 22138 16164 22172
rect 16102 22104 16118 22138
rect 16152 22104 16164 22138
rect 16102 22070 16164 22104
rect 16102 22036 16118 22070
rect 16152 22036 16164 22070
rect 16102 22002 16164 22036
rect 16102 21968 16118 22002
rect 16152 21968 16164 22002
rect 16102 21934 16164 21968
rect 16102 21900 16118 21934
rect 16152 21900 16164 21934
rect 16102 21866 16164 21900
rect 16102 21832 16118 21866
rect 16152 21832 16164 21866
rect 16102 21798 16164 21832
rect 16102 21764 16118 21798
rect 16152 21764 16164 21798
rect 16102 21730 16164 21764
rect 16102 21696 16118 21730
rect 16152 21696 16164 21730
rect 16102 21662 16164 21696
rect 16102 21628 16118 21662
rect 16152 21628 16164 21662
rect 16102 21594 16164 21628
rect 16102 21560 16118 21594
rect 16152 21560 16164 21594
rect 16102 21526 16164 21560
rect 16102 21492 16118 21526
rect 16152 21492 16164 21526
rect 16102 21458 16164 21492
rect 16102 21424 16118 21458
rect 16152 21424 16164 21458
rect 16102 21390 16164 21424
rect 16102 21356 16118 21390
rect 16152 21356 16164 21390
rect 16102 21322 16164 21356
rect 16102 21288 16118 21322
rect 16152 21288 16164 21322
rect 16102 21254 16164 21288
rect 16102 21220 16118 21254
rect 16152 21220 16164 21254
rect 16102 21189 16164 21220
rect 17080 15912 17142 15943
rect 17080 15878 17092 15912
rect 17126 15878 17142 15912
rect 17080 15844 17142 15878
rect 17080 15810 17092 15844
rect 17126 15810 17142 15844
rect 17080 15776 17142 15810
rect 17080 15742 17092 15776
rect 17126 15742 17142 15776
rect 17080 15708 17142 15742
rect 17080 15674 17092 15708
rect 17126 15674 17142 15708
rect 17080 15640 17142 15674
rect 17080 15606 17092 15640
rect 17126 15606 17142 15640
rect 17080 15572 17142 15606
rect 17080 15538 17092 15572
rect 17126 15538 17142 15572
rect 17080 15504 17142 15538
rect 17080 15470 17092 15504
rect 17126 15470 17142 15504
rect 17080 15436 17142 15470
rect 17080 15402 17092 15436
rect 17126 15402 17142 15436
rect 17080 15368 17142 15402
rect 17080 15334 17092 15368
rect 17126 15334 17142 15368
rect 17080 15300 17142 15334
rect 17080 15266 17092 15300
rect 17126 15266 17142 15300
rect 17080 15232 17142 15266
rect 17080 15198 17092 15232
rect 17126 15198 17142 15232
rect 17080 15164 17142 15198
rect 17080 15130 17092 15164
rect 17126 15130 17142 15164
rect 17080 15096 17142 15130
rect 17080 15062 17092 15096
rect 17126 15062 17142 15096
rect 17080 15028 17142 15062
rect 17080 14994 17092 15028
rect 17126 14994 17142 15028
rect 17080 14960 17142 14994
rect 17080 14926 17092 14960
rect 17126 14926 17142 14960
rect 17080 14892 17142 14926
rect 17080 14858 17092 14892
rect 17126 14858 17142 14892
rect 17080 14824 17142 14858
rect 17080 14790 17092 14824
rect 17126 14790 17142 14824
rect 17080 14756 17142 14790
rect 17080 14722 17092 14756
rect 17126 14722 17142 14756
rect 17080 14688 17142 14722
rect 17080 14654 17092 14688
rect 17126 14654 17142 14688
rect 17080 14620 17142 14654
rect 17080 14586 17092 14620
rect 17126 14586 17142 14620
rect 17080 14552 17142 14586
rect 17080 14518 17092 14552
rect 17126 14518 17142 14552
rect 17080 14484 17142 14518
rect 17080 14450 17092 14484
rect 17126 14450 17142 14484
rect 17080 14416 17142 14450
rect 17080 14382 17092 14416
rect 17126 14382 17142 14416
rect 17080 14348 17142 14382
rect 17080 14314 17092 14348
rect 17126 14314 17142 14348
rect 17080 14280 17142 14314
rect 17080 14246 17092 14280
rect 17126 14246 17142 14280
rect 17080 14212 17142 14246
rect 17080 14178 17092 14212
rect 17126 14178 17142 14212
rect 17080 14144 17142 14178
rect 17080 14110 17092 14144
rect 17126 14110 17142 14144
rect 17080 14076 17142 14110
rect 17080 14042 17092 14076
rect 17126 14042 17142 14076
rect 17080 14008 17142 14042
rect 17080 13974 17092 14008
rect 17126 13974 17142 14008
rect 17080 13943 17142 13974
rect 17172 15912 17238 15943
rect 17172 15878 17188 15912
rect 17222 15878 17238 15912
rect 17172 15844 17238 15878
rect 17172 15810 17188 15844
rect 17222 15810 17238 15844
rect 17172 15776 17238 15810
rect 17172 15742 17188 15776
rect 17222 15742 17238 15776
rect 17172 15708 17238 15742
rect 17172 15674 17188 15708
rect 17222 15674 17238 15708
rect 17172 15640 17238 15674
rect 17172 15606 17188 15640
rect 17222 15606 17238 15640
rect 17172 15572 17238 15606
rect 17172 15538 17188 15572
rect 17222 15538 17238 15572
rect 17172 15504 17238 15538
rect 17172 15470 17188 15504
rect 17222 15470 17238 15504
rect 17172 15436 17238 15470
rect 17172 15402 17188 15436
rect 17222 15402 17238 15436
rect 17172 15368 17238 15402
rect 17172 15334 17188 15368
rect 17222 15334 17238 15368
rect 17172 15300 17238 15334
rect 17172 15266 17188 15300
rect 17222 15266 17238 15300
rect 17172 15232 17238 15266
rect 17172 15198 17188 15232
rect 17222 15198 17238 15232
rect 17172 15164 17238 15198
rect 17172 15130 17188 15164
rect 17222 15130 17238 15164
rect 17172 15096 17238 15130
rect 17172 15062 17188 15096
rect 17222 15062 17238 15096
rect 17172 15028 17238 15062
rect 17172 14994 17188 15028
rect 17222 14994 17238 15028
rect 17172 14960 17238 14994
rect 17172 14926 17188 14960
rect 17222 14926 17238 14960
rect 17172 14892 17238 14926
rect 17172 14858 17188 14892
rect 17222 14858 17238 14892
rect 17172 14824 17238 14858
rect 17172 14790 17188 14824
rect 17222 14790 17238 14824
rect 17172 14756 17238 14790
rect 17172 14722 17188 14756
rect 17222 14722 17238 14756
rect 17172 14688 17238 14722
rect 17172 14654 17188 14688
rect 17222 14654 17238 14688
rect 17172 14620 17238 14654
rect 17172 14586 17188 14620
rect 17222 14586 17238 14620
rect 17172 14552 17238 14586
rect 17172 14518 17188 14552
rect 17222 14518 17238 14552
rect 17172 14484 17238 14518
rect 17172 14450 17188 14484
rect 17222 14450 17238 14484
rect 17172 14416 17238 14450
rect 17172 14382 17188 14416
rect 17222 14382 17238 14416
rect 17172 14348 17238 14382
rect 17172 14314 17188 14348
rect 17222 14314 17238 14348
rect 17172 14280 17238 14314
rect 17172 14246 17188 14280
rect 17222 14246 17238 14280
rect 17172 14212 17238 14246
rect 17172 14178 17188 14212
rect 17222 14178 17238 14212
rect 17172 14144 17238 14178
rect 17172 14110 17188 14144
rect 17222 14110 17238 14144
rect 17172 14076 17238 14110
rect 17172 14042 17188 14076
rect 17222 14042 17238 14076
rect 17172 14008 17238 14042
rect 17172 13974 17188 14008
rect 17222 13974 17238 14008
rect 17172 13943 17238 13974
rect 17268 15912 17334 15943
rect 17268 15878 17284 15912
rect 17318 15878 17334 15912
rect 17268 15844 17334 15878
rect 17268 15810 17284 15844
rect 17318 15810 17334 15844
rect 17268 15776 17334 15810
rect 17268 15742 17284 15776
rect 17318 15742 17334 15776
rect 17268 15708 17334 15742
rect 17268 15674 17284 15708
rect 17318 15674 17334 15708
rect 17268 15640 17334 15674
rect 17268 15606 17284 15640
rect 17318 15606 17334 15640
rect 17268 15572 17334 15606
rect 17268 15538 17284 15572
rect 17318 15538 17334 15572
rect 17268 15504 17334 15538
rect 17268 15470 17284 15504
rect 17318 15470 17334 15504
rect 17268 15436 17334 15470
rect 17268 15402 17284 15436
rect 17318 15402 17334 15436
rect 17268 15368 17334 15402
rect 17268 15334 17284 15368
rect 17318 15334 17334 15368
rect 17268 15300 17334 15334
rect 17268 15266 17284 15300
rect 17318 15266 17334 15300
rect 17268 15232 17334 15266
rect 17268 15198 17284 15232
rect 17318 15198 17334 15232
rect 17268 15164 17334 15198
rect 17268 15130 17284 15164
rect 17318 15130 17334 15164
rect 17268 15096 17334 15130
rect 17268 15062 17284 15096
rect 17318 15062 17334 15096
rect 17268 15028 17334 15062
rect 17268 14994 17284 15028
rect 17318 14994 17334 15028
rect 17268 14960 17334 14994
rect 17268 14926 17284 14960
rect 17318 14926 17334 14960
rect 17268 14892 17334 14926
rect 17268 14858 17284 14892
rect 17318 14858 17334 14892
rect 17268 14824 17334 14858
rect 17268 14790 17284 14824
rect 17318 14790 17334 14824
rect 17268 14756 17334 14790
rect 17268 14722 17284 14756
rect 17318 14722 17334 14756
rect 17268 14688 17334 14722
rect 17268 14654 17284 14688
rect 17318 14654 17334 14688
rect 17268 14620 17334 14654
rect 17268 14586 17284 14620
rect 17318 14586 17334 14620
rect 17268 14552 17334 14586
rect 17268 14518 17284 14552
rect 17318 14518 17334 14552
rect 17268 14484 17334 14518
rect 17268 14450 17284 14484
rect 17318 14450 17334 14484
rect 17268 14416 17334 14450
rect 17268 14382 17284 14416
rect 17318 14382 17334 14416
rect 17268 14348 17334 14382
rect 17268 14314 17284 14348
rect 17318 14314 17334 14348
rect 17268 14280 17334 14314
rect 17268 14246 17284 14280
rect 17318 14246 17334 14280
rect 17268 14212 17334 14246
rect 17268 14178 17284 14212
rect 17318 14178 17334 14212
rect 17268 14144 17334 14178
rect 17268 14110 17284 14144
rect 17318 14110 17334 14144
rect 17268 14076 17334 14110
rect 17268 14042 17284 14076
rect 17318 14042 17334 14076
rect 17268 14008 17334 14042
rect 17268 13974 17284 14008
rect 17318 13974 17334 14008
rect 17268 13943 17334 13974
rect 17364 15912 17426 15943
rect 17364 15878 17380 15912
rect 17414 15878 17426 15912
rect 17364 15844 17426 15878
rect 17364 15810 17380 15844
rect 17414 15810 17426 15844
rect 17364 15776 17426 15810
rect 17364 15742 17380 15776
rect 17414 15742 17426 15776
rect 17364 15708 17426 15742
rect 17364 15674 17380 15708
rect 17414 15674 17426 15708
rect 17364 15640 17426 15674
rect 17364 15606 17380 15640
rect 17414 15606 17426 15640
rect 17364 15572 17426 15606
rect 17364 15538 17380 15572
rect 17414 15538 17426 15572
rect 17364 15504 17426 15538
rect 17364 15470 17380 15504
rect 17414 15470 17426 15504
rect 17364 15436 17426 15470
rect 17364 15402 17380 15436
rect 17414 15402 17426 15436
rect 17364 15368 17426 15402
rect 17364 15334 17380 15368
rect 17414 15334 17426 15368
rect 17364 15300 17426 15334
rect 17364 15266 17380 15300
rect 17414 15266 17426 15300
rect 17364 15232 17426 15266
rect 17364 15198 17380 15232
rect 17414 15198 17426 15232
rect 17364 15164 17426 15198
rect 17364 15130 17380 15164
rect 17414 15130 17426 15164
rect 17364 15096 17426 15130
rect 17364 15062 17380 15096
rect 17414 15062 17426 15096
rect 17364 15028 17426 15062
rect 17364 14994 17380 15028
rect 17414 14994 17426 15028
rect 17364 14960 17426 14994
rect 17364 14926 17380 14960
rect 17414 14926 17426 14960
rect 17364 14892 17426 14926
rect 17364 14858 17380 14892
rect 17414 14858 17426 14892
rect 17364 14824 17426 14858
rect 17364 14790 17380 14824
rect 17414 14790 17426 14824
rect 17364 14756 17426 14790
rect 17364 14722 17380 14756
rect 17414 14722 17426 14756
rect 17364 14688 17426 14722
rect 17364 14654 17380 14688
rect 17414 14654 17426 14688
rect 17364 14620 17426 14654
rect 17364 14586 17380 14620
rect 17414 14586 17426 14620
rect 17364 14552 17426 14586
rect 17364 14518 17380 14552
rect 17414 14518 17426 14552
rect 17364 14484 17426 14518
rect 17364 14450 17380 14484
rect 17414 14450 17426 14484
rect 17364 14416 17426 14450
rect 17364 14382 17380 14416
rect 17414 14382 17426 14416
rect 17364 14348 17426 14382
rect 17364 14314 17380 14348
rect 17414 14314 17426 14348
rect 17364 14280 17426 14314
rect 17364 14246 17380 14280
rect 17414 14246 17426 14280
rect 17364 14212 17426 14246
rect 17364 14178 17380 14212
rect 17414 14178 17426 14212
rect 17364 14144 17426 14178
rect 17364 14110 17380 14144
rect 17414 14110 17426 14144
rect 17364 14076 17426 14110
rect 17364 14042 17380 14076
rect 17414 14042 17426 14076
rect 17364 14008 17426 14042
rect 17364 13974 17380 14008
rect 17414 13974 17426 14008
rect 17364 13943 17426 13974
<< ndiffc >>
rect 13970 23085 14004 23119
rect 13970 23017 14004 23051
rect 13970 22949 14004 22983
rect 13970 22881 14004 22915
rect 13970 22813 14004 22847
rect 13970 22745 14004 22779
rect 13970 22677 14004 22711
rect 13970 22609 14004 22643
rect 13970 22541 14004 22575
rect 13970 22473 14004 22507
rect 13970 22405 14004 22439
rect 13970 22337 14004 22371
rect 13970 22269 14004 22303
rect 13970 22201 14004 22235
rect 13970 22133 14004 22167
rect 13970 22065 14004 22099
rect 13970 21997 14004 22031
rect 13970 21929 14004 21963
rect 13970 21861 14004 21895
rect 13970 21793 14004 21827
rect 13970 21725 14004 21759
rect 13970 21657 14004 21691
rect 13970 21589 14004 21623
rect 13970 21521 14004 21555
rect 13970 21453 14004 21487
rect 13970 21385 14004 21419
rect 13970 21317 14004 21351
rect 13970 21249 14004 21283
rect 13970 21181 14004 21215
rect 14066 23085 14100 23119
rect 14066 23017 14100 23051
rect 14066 22949 14100 22983
rect 14066 22881 14100 22915
rect 14066 22813 14100 22847
rect 14066 22745 14100 22779
rect 14066 22677 14100 22711
rect 14066 22609 14100 22643
rect 14066 22541 14100 22575
rect 14066 22473 14100 22507
rect 14066 22405 14100 22439
rect 14066 22337 14100 22371
rect 14066 22269 14100 22303
rect 14066 22201 14100 22235
rect 14066 22133 14100 22167
rect 14066 22065 14100 22099
rect 14066 21997 14100 22031
rect 14066 21929 14100 21963
rect 14066 21861 14100 21895
rect 14066 21793 14100 21827
rect 14066 21725 14100 21759
rect 14066 21657 14100 21691
rect 14066 21589 14100 21623
rect 14066 21521 14100 21555
rect 14066 21453 14100 21487
rect 14066 21385 14100 21419
rect 14066 21317 14100 21351
rect 14066 21249 14100 21283
rect 14066 21181 14100 21215
rect 14162 23085 14196 23119
rect 14162 23017 14196 23051
rect 14162 22949 14196 22983
rect 14162 22881 14196 22915
rect 14162 22813 14196 22847
rect 14162 22745 14196 22779
rect 14162 22677 14196 22711
rect 14162 22609 14196 22643
rect 14162 22541 14196 22575
rect 14162 22473 14196 22507
rect 14162 22405 14196 22439
rect 14162 22337 14196 22371
rect 14162 22269 14196 22303
rect 14162 22201 14196 22235
rect 14162 22133 14196 22167
rect 14162 22065 14196 22099
rect 14162 21997 14196 22031
rect 14162 21929 14196 21963
rect 14162 21861 14196 21895
rect 14162 21793 14196 21827
rect 14162 21725 14196 21759
rect 14162 21657 14196 21691
rect 14162 21589 14196 21623
rect 14162 21521 14196 21555
rect 14162 21453 14196 21487
rect 14162 21385 14196 21419
rect 14162 21317 14196 21351
rect 14162 21249 14196 21283
rect 14162 21181 14196 21215
rect 14258 23085 14292 23119
rect 14258 23017 14292 23051
rect 14258 22949 14292 22983
rect 14258 22881 14292 22915
rect 14258 22813 14292 22847
rect 14258 22745 14292 22779
rect 14258 22677 14292 22711
rect 14258 22609 14292 22643
rect 14258 22541 14292 22575
rect 14258 22473 14292 22507
rect 14258 22405 14292 22439
rect 14258 22337 14292 22371
rect 14258 22269 14292 22303
rect 14258 22201 14292 22235
rect 14258 22133 14292 22167
rect 14258 22065 14292 22099
rect 14258 21997 14292 22031
rect 14258 21929 14292 21963
rect 14258 21861 14292 21895
rect 14258 21793 14292 21827
rect 14258 21725 14292 21759
rect 14258 21657 14292 21691
rect 14258 21589 14292 21623
rect 14258 21521 14292 21555
rect 14258 21453 14292 21487
rect 14258 21385 14292 21419
rect 14258 21317 14292 21351
rect 14258 21249 14292 21283
rect 14258 21181 14292 21215
rect 14354 23085 14388 23119
rect 14354 23017 14388 23051
rect 14354 22949 14388 22983
rect 14354 22881 14388 22915
rect 14354 22813 14388 22847
rect 14354 22745 14388 22779
rect 14354 22677 14388 22711
rect 14354 22609 14388 22643
rect 14354 22541 14388 22575
rect 14354 22473 14388 22507
rect 14354 22405 14388 22439
rect 14354 22337 14388 22371
rect 14354 22269 14388 22303
rect 14354 22201 14388 22235
rect 14354 22133 14388 22167
rect 14354 22065 14388 22099
rect 14354 21997 14388 22031
rect 14354 21929 14388 21963
rect 14354 21861 14388 21895
rect 14354 21793 14388 21827
rect 14354 21725 14388 21759
rect 14354 21657 14388 21691
rect 14354 21589 14388 21623
rect 14354 21521 14388 21555
rect 14354 21453 14388 21487
rect 14354 21385 14388 21419
rect 14354 21317 14388 21351
rect 14354 21249 14388 21283
rect 14354 21181 14388 21215
rect 14450 23085 14484 23119
rect 14450 23017 14484 23051
rect 14450 22949 14484 22983
rect 14450 22881 14484 22915
rect 14450 22813 14484 22847
rect 14450 22745 14484 22779
rect 14450 22677 14484 22711
rect 14450 22609 14484 22643
rect 14450 22541 14484 22575
rect 14450 22473 14484 22507
rect 14450 22405 14484 22439
rect 14450 22337 14484 22371
rect 14450 22269 14484 22303
rect 14450 22201 14484 22235
rect 14450 22133 14484 22167
rect 14450 22065 14484 22099
rect 14450 21997 14484 22031
rect 14450 21929 14484 21963
rect 14450 21861 14484 21895
rect 14450 21793 14484 21827
rect 14450 21725 14484 21759
rect 14450 21657 14484 21691
rect 14450 21589 14484 21623
rect 14450 21521 14484 21555
rect 14450 21453 14484 21487
rect 14450 21385 14484 21419
rect 14450 21317 14484 21351
rect 14450 21249 14484 21283
rect 14450 21181 14484 21215
rect 14546 23085 14580 23119
rect 14546 23017 14580 23051
rect 14546 22949 14580 22983
rect 14546 22881 14580 22915
rect 14546 22813 14580 22847
rect 14546 22745 14580 22779
rect 14546 22677 14580 22711
rect 14546 22609 14580 22643
rect 14546 22541 14580 22575
rect 14546 22473 14580 22507
rect 14546 22405 14580 22439
rect 14546 22337 14580 22371
rect 14546 22269 14580 22303
rect 14546 22201 14580 22235
rect 14546 22133 14580 22167
rect 14546 22065 14580 22099
rect 14546 21997 14580 22031
rect 14546 21929 14580 21963
rect 14546 21861 14580 21895
rect 14546 21793 14580 21827
rect 14546 21725 14580 21759
rect 14546 21657 14580 21691
rect 14546 21589 14580 21623
rect 14546 21521 14580 21555
rect 14546 21453 14580 21487
rect 14546 21385 14580 21419
rect 14546 21317 14580 21351
rect 14546 21249 14580 21283
rect 14546 21181 14580 21215
rect 14642 23085 14676 23119
rect 14642 23017 14676 23051
rect 14642 22949 14676 22983
rect 14642 22881 14676 22915
rect 14642 22813 14676 22847
rect 14642 22745 14676 22779
rect 14642 22677 14676 22711
rect 14642 22609 14676 22643
rect 14642 22541 14676 22575
rect 14642 22473 14676 22507
rect 14642 22405 14676 22439
rect 14642 22337 14676 22371
rect 14642 22269 14676 22303
rect 14642 22201 14676 22235
rect 14642 22133 14676 22167
rect 14642 22065 14676 22099
rect 14642 21997 14676 22031
rect 14642 21929 14676 21963
rect 14642 21861 14676 21895
rect 14642 21793 14676 21827
rect 14642 21725 14676 21759
rect 14642 21657 14676 21691
rect 14642 21589 14676 21623
rect 14642 21521 14676 21555
rect 14642 21453 14676 21487
rect 14642 21385 14676 21419
rect 14642 21317 14676 21351
rect 14642 21249 14676 21283
rect 14642 21181 14676 21215
rect 14738 23085 14772 23119
rect 14738 23017 14772 23051
rect 14738 22949 14772 22983
rect 14738 22881 14772 22915
rect 14738 22813 14772 22847
rect 14738 22745 14772 22779
rect 14738 22677 14772 22711
rect 14738 22609 14772 22643
rect 14738 22541 14772 22575
rect 14738 22473 14772 22507
rect 14738 22405 14772 22439
rect 14738 22337 14772 22371
rect 14738 22269 14772 22303
rect 14738 22201 14772 22235
rect 14738 22133 14772 22167
rect 14738 22065 14772 22099
rect 14738 21997 14772 22031
rect 14738 21929 14772 21963
rect 14738 21861 14772 21895
rect 14738 21793 14772 21827
rect 14738 21725 14772 21759
rect 14738 21657 14772 21691
rect 14738 21589 14772 21623
rect 14738 21521 14772 21555
rect 14738 21453 14772 21487
rect 14738 21385 14772 21419
rect 14738 21317 14772 21351
rect 14738 21249 14772 21283
rect 14738 21181 14772 21215
rect 16662 23975 16696 24009
rect 16662 23907 16696 23941
rect 16662 23839 16696 23873
rect 16662 23771 16696 23805
rect 16662 23703 16696 23737
rect 16662 23635 16696 23669
rect 16662 23567 16696 23601
rect 16662 23499 16696 23533
rect 16662 23431 16696 23465
rect 16662 23363 16696 23397
rect 16662 23295 16696 23329
rect 16662 23227 16696 23261
rect 16662 23159 16696 23193
rect 16662 23091 16696 23125
rect 16662 23023 16696 23057
rect 16662 22955 16696 22989
rect 16662 22887 16696 22921
rect 16662 22819 16696 22853
rect 16662 22751 16696 22785
rect 16662 22683 16696 22717
rect 16662 22615 16696 22649
rect 16662 22547 16696 22581
rect 16662 22479 16696 22513
rect 16662 22411 16696 22445
rect 16662 22343 16696 22377
rect 16662 22275 16696 22309
rect 16662 22207 16696 22241
rect 16662 22139 16696 22173
rect 16662 22071 16696 22105
rect 16758 23975 16792 24009
rect 16758 23907 16792 23941
rect 16758 23839 16792 23873
rect 16758 23771 16792 23805
rect 16758 23703 16792 23737
rect 16758 23635 16792 23669
rect 16758 23567 16792 23601
rect 16758 23499 16792 23533
rect 16758 23431 16792 23465
rect 16758 23363 16792 23397
rect 16758 23295 16792 23329
rect 16758 23227 16792 23261
rect 16758 23159 16792 23193
rect 16758 23091 16792 23125
rect 16758 23023 16792 23057
rect 16758 22955 16792 22989
rect 16758 22887 16792 22921
rect 16758 22819 16792 22853
rect 16758 22751 16792 22785
rect 16758 22683 16792 22717
rect 16758 22615 16792 22649
rect 16758 22547 16792 22581
rect 16758 22479 16792 22513
rect 16758 22411 16792 22445
rect 16758 22343 16792 22377
rect 16758 22275 16792 22309
rect 16758 22207 16792 22241
rect 16758 22139 16792 22173
rect 16758 22071 16792 22105
rect 16854 23975 16888 24009
rect 16854 23907 16888 23941
rect 16854 23839 16888 23873
rect 16854 23771 16888 23805
rect 16854 23703 16888 23737
rect 16854 23635 16888 23669
rect 16854 23567 16888 23601
rect 16854 23499 16888 23533
rect 16854 23431 16888 23465
rect 16854 23363 16888 23397
rect 16854 23295 16888 23329
rect 16854 23227 16888 23261
rect 16854 23159 16888 23193
rect 16854 23091 16888 23125
rect 16854 23023 16888 23057
rect 16854 22955 16888 22989
rect 16854 22887 16888 22921
rect 16854 22819 16888 22853
rect 16854 22751 16888 22785
rect 16854 22683 16888 22717
rect 16854 22615 16888 22649
rect 16854 22547 16888 22581
rect 16854 22479 16888 22513
rect 16854 22411 16888 22445
rect 16854 22343 16888 22377
rect 16854 22275 16888 22309
rect 16854 22207 16888 22241
rect 16854 22139 16888 22173
rect 16854 22071 16888 22105
rect 16950 23975 16984 24009
rect 16950 23907 16984 23941
rect 16950 23839 16984 23873
rect 16950 23771 16984 23805
rect 16950 23703 16984 23737
rect 16950 23635 16984 23669
rect 16950 23567 16984 23601
rect 16950 23499 16984 23533
rect 16950 23431 16984 23465
rect 16950 23363 16984 23397
rect 16950 23295 16984 23329
rect 16950 23227 16984 23261
rect 16950 23159 16984 23193
rect 16950 23091 16984 23125
rect 16950 23023 16984 23057
rect 16950 22955 16984 22989
rect 16950 22887 16984 22921
rect 16950 22819 16984 22853
rect 16950 22751 16984 22785
rect 16950 22683 16984 22717
rect 16950 22615 16984 22649
rect 16950 22547 16984 22581
rect 16950 22479 16984 22513
rect 16950 22411 16984 22445
rect 16950 22343 16984 22377
rect 16950 22275 16984 22309
rect 16950 22207 16984 22241
rect 16950 22139 16984 22173
rect 16950 22071 16984 22105
rect 17046 23975 17080 24009
rect 17046 23907 17080 23941
rect 17046 23839 17080 23873
rect 17046 23771 17080 23805
rect 17046 23703 17080 23737
rect 17046 23635 17080 23669
rect 17046 23567 17080 23601
rect 17046 23499 17080 23533
rect 17046 23431 17080 23465
rect 17046 23363 17080 23397
rect 17046 23295 17080 23329
rect 17046 23227 17080 23261
rect 17046 23159 17080 23193
rect 17046 23091 17080 23125
rect 17046 23023 17080 23057
rect 17046 22955 17080 22989
rect 17046 22887 17080 22921
rect 17046 22819 17080 22853
rect 17046 22751 17080 22785
rect 17046 22683 17080 22717
rect 17046 22615 17080 22649
rect 17046 22547 17080 22581
rect 17046 22479 17080 22513
rect 17046 22411 17080 22445
rect 17046 22343 17080 22377
rect 17046 22275 17080 22309
rect 17046 22207 17080 22241
rect 17046 22139 17080 22173
rect 17046 22071 17080 22105
rect 17142 23975 17176 24009
rect 17142 23907 17176 23941
rect 17142 23839 17176 23873
rect 17142 23771 17176 23805
rect 17142 23703 17176 23737
rect 17142 23635 17176 23669
rect 17142 23567 17176 23601
rect 17142 23499 17176 23533
rect 17142 23431 17176 23465
rect 17142 23363 17176 23397
rect 17142 23295 17176 23329
rect 17142 23227 17176 23261
rect 17142 23159 17176 23193
rect 17142 23091 17176 23125
rect 17142 23023 17176 23057
rect 17142 22955 17176 22989
rect 17142 22887 17176 22921
rect 17142 22819 17176 22853
rect 17142 22751 17176 22785
rect 17142 22683 17176 22717
rect 17142 22615 17176 22649
rect 17142 22547 17176 22581
rect 17142 22479 17176 22513
rect 17142 22411 17176 22445
rect 17142 22343 17176 22377
rect 17142 22275 17176 22309
rect 17142 22207 17176 22241
rect 17142 22139 17176 22173
rect 17142 22071 17176 22105
rect 17238 23975 17272 24009
rect 17238 23907 17272 23941
rect 17238 23839 17272 23873
rect 17238 23771 17272 23805
rect 17238 23703 17272 23737
rect 17238 23635 17272 23669
rect 17238 23567 17272 23601
rect 17238 23499 17272 23533
rect 17238 23431 17272 23465
rect 17238 23363 17272 23397
rect 17238 23295 17272 23329
rect 17238 23227 17272 23261
rect 17238 23159 17272 23193
rect 17238 23091 17272 23125
rect 17238 23023 17272 23057
rect 17238 22955 17272 22989
rect 17238 22887 17272 22921
rect 17238 22819 17272 22853
rect 17238 22751 17272 22785
rect 17238 22683 17272 22717
rect 17238 22615 17272 22649
rect 17238 22547 17272 22581
rect 17238 22479 17272 22513
rect 17238 22411 17272 22445
rect 17238 22343 17272 22377
rect 17238 22275 17272 22309
rect 17238 22207 17272 22241
rect 17238 22139 17272 22173
rect 17238 22071 17272 22105
rect 17334 23975 17368 24009
rect 17334 23907 17368 23941
rect 17334 23839 17368 23873
rect 17334 23771 17368 23805
rect 17334 23703 17368 23737
rect 17334 23635 17368 23669
rect 17334 23567 17368 23601
rect 17334 23499 17368 23533
rect 17334 23431 17368 23465
rect 17334 23363 17368 23397
rect 17334 23295 17368 23329
rect 17334 23227 17368 23261
rect 17334 23159 17368 23193
rect 17334 23091 17368 23125
rect 17334 23023 17368 23057
rect 17334 22955 17368 22989
rect 17334 22887 17368 22921
rect 17334 22819 17368 22853
rect 17334 22751 17368 22785
rect 17334 22683 17368 22717
rect 17334 22615 17368 22649
rect 17334 22547 17368 22581
rect 17334 22479 17368 22513
rect 17334 22411 17368 22445
rect 17334 22343 17368 22377
rect 17334 22275 17368 22309
rect 17334 22207 17368 22241
rect 17334 22139 17368 22173
rect 17334 22071 17368 22105
rect 17430 23975 17464 24009
rect 17430 23907 17464 23941
rect 17430 23839 17464 23873
rect 17430 23771 17464 23805
rect 17430 23703 17464 23737
rect 17430 23635 17464 23669
rect 17430 23567 17464 23601
rect 17430 23499 17464 23533
rect 17430 23431 17464 23465
rect 17430 23363 17464 23397
rect 17430 23295 17464 23329
rect 17430 23227 17464 23261
rect 17430 23159 17464 23193
rect 17430 23091 17464 23125
rect 17430 23023 17464 23057
rect 17430 22955 17464 22989
rect 17430 22887 17464 22921
rect 17430 22819 17464 22853
rect 17430 22751 17464 22785
rect 17430 22683 17464 22717
rect 17430 22615 17464 22649
rect 17430 22547 17464 22581
rect 17430 22479 17464 22513
rect 17430 22411 17464 22445
rect 17430 22343 17464 22377
rect 17430 22275 17464 22309
rect 17430 22207 17464 22241
rect 17430 22139 17464 22173
rect 17430 22071 17464 22105
rect 17526 23975 17560 24009
rect 17526 23907 17560 23941
rect 17526 23839 17560 23873
rect 17526 23771 17560 23805
rect 17526 23703 17560 23737
rect 17526 23635 17560 23669
rect 17526 23567 17560 23601
rect 17526 23499 17560 23533
rect 17526 23431 17560 23465
rect 17526 23363 17560 23397
rect 17526 23295 17560 23329
rect 17526 23227 17560 23261
rect 17526 23159 17560 23193
rect 17526 23091 17560 23125
rect 17526 23023 17560 23057
rect 17526 22955 17560 22989
rect 17526 22887 17560 22921
rect 17526 22819 17560 22853
rect 17526 22751 17560 22785
rect 17526 22683 17560 22717
rect 17526 22615 17560 22649
rect 17526 22547 17560 22581
rect 17526 22479 17560 22513
rect 17526 22411 17560 22445
rect 17526 22343 17560 22377
rect 17526 22275 17560 22309
rect 17526 22207 17560 22241
rect 17526 22139 17560 22173
rect 17526 22071 17560 22105
rect 17622 23975 17656 24009
rect 17622 23907 17656 23941
rect 17622 23839 17656 23873
rect 17622 23771 17656 23805
rect 17622 23703 17656 23737
rect 17622 23635 17656 23669
rect 17622 23567 17656 23601
rect 17622 23499 17656 23533
rect 17622 23431 17656 23465
rect 17622 23363 17656 23397
rect 17622 23295 17656 23329
rect 17622 23227 17656 23261
rect 17622 23159 17656 23193
rect 17622 23091 17656 23125
rect 17622 23023 17656 23057
rect 17622 22955 17656 22989
rect 17622 22887 17656 22921
rect 17622 22819 17656 22853
rect 17622 22751 17656 22785
rect 17622 22683 17656 22717
rect 17622 22615 17656 22649
rect 17622 22547 17656 22581
rect 17622 22479 17656 22513
rect 17622 22411 17656 22445
rect 17622 22343 17656 22377
rect 17622 22275 17656 22309
rect 17622 22207 17656 22241
rect 17622 22139 17656 22173
rect 17622 22071 17656 22105
rect 14830 20398 14864 20432
rect 14830 20330 14864 20364
rect 14830 20262 14864 20296
rect 14830 20194 14864 20228
rect 14830 20126 14864 20160
rect 14830 20058 14864 20092
rect 14830 19990 14864 20024
rect 14830 19922 14864 19956
rect 14830 19854 14864 19888
rect 14830 19786 14864 19820
rect 14830 19718 14864 19752
rect 14830 19650 14864 19684
rect 14830 19582 14864 19616
rect 14830 19514 14864 19548
rect 14830 19446 14864 19480
rect 14830 19378 14864 19412
rect 14830 19310 14864 19344
rect 14830 19242 14864 19276
rect 14830 19174 14864 19208
rect 14926 20398 14960 20432
rect 14926 20330 14960 20364
rect 14926 20262 14960 20296
rect 14926 20194 14960 20228
rect 14926 20126 14960 20160
rect 14926 20058 14960 20092
rect 14926 19990 14960 20024
rect 14926 19922 14960 19956
rect 14926 19854 14960 19888
rect 14926 19786 14960 19820
rect 14926 19718 14960 19752
rect 14926 19650 14960 19684
rect 14926 19582 14960 19616
rect 14926 19514 14960 19548
rect 14926 19446 14960 19480
rect 14926 19378 14960 19412
rect 14926 19310 14960 19344
rect 14926 19242 14960 19276
rect 14926 19174 14960 19208
rect 15022 20398 15056 20432
rect 15022 20330 15056 20364
rect 15022 20262 15056 20296
rect 15022 20194 15056 20228
rect 15022 20126 15056 20160
rect 15022 20058 15056 20092
rect 15022 19990 15056 20024
rect 15022 19922 15056 19956
rect 15022 19854 15056 19888
rect 15022 19786 15056 19820
rect 15022 19718 15056 19752
rect 15022 19650 15056 19684
rect 15022 19582 15056 19616
rect 15022 19514 15056 19548
rect 15022 19446 15056 19480
rect 15022 19378 15056 19412
rect 15022 19310 15056 19344
rect 15022 19242 15056 19276
rect 15022 19174 15056 19208
rect 15118 20398 15152 20432
rect 15118 20330 15152 20364
rect 15118 20262 15152 20296
rect 15118 20194 15152 20228
rect 15118 20126 15152 20160
rect 15118 20058 15152 20092
rect 15118 19990 15152 20024
rect 15118 19922 15152 19956
rect 15118 19854 15152 19888
rect 15118 19786 15152 19820
rect 15118 19718 15152 19752
rect 15118 19650 15152 19684
rect 15118 19582 15152 19616
rect 15118 19514 15152 19548
rect 15118 19446 15152 19480
rect 15118 19378 15152 19412
rect 15118 19310 15152 19344
rect 15118 19242 15152 19276
rect 15118 19174 15152 19208
rect 15214 20398 15248 20432
rect 15214 20330 15248 20364
rect 15214 20262 15248 20296
rect 15214 20194 15248 20228
rect 15214 20126 15248 20160
rect 15214 20058 15248 20092
rect 15214 19990 15248 20024
rect 15214 19922 15248 19956
rect 15214 19854 15248 19888
rect 15214 19786 15248 19820
rect 15214 19718 15248 19752
rect 15214 19650 15248 19684
rect 15214 19582 15248 19616
rect 15214 19514 15248 19548
rect 15214 19446 15248 19480
rect 15214 19378 15248 19412
rect 15214 19310 15248 19344
rect 15214 19242 15248 19276
rect 15214 19174 15248 19208
rect 15310 20398 15344 20432
rect 15310 20330 15344 20364
rect 15310 20262 15344 20296
rect 15310 20194 15344 20228
rect 15310 20126 15344 20160
rect 15310 20058 15344 20092
rect 15310 19990 15344 20024
rect 15310 19922 15344 19956
rect 15310 19854 15344 19888
rect 15310 19786 15344 19820
rect 15310 19718 15344 19752
rect 15310 19650 15344 19684
rect 15310 19582 15344 19616
rect 15310 19514 15344 19548
rect 15310 19446 15344 19480
rect 15310 19378 15344 19412
rect 15310 19310 15344 19344
rect 15310 19242 15344 19276
rect 15310 19174 15344 19208
rect 15406 20398 15440 20432
rect 15406 20330 15440 20364
rect 15406 20262 15440 20296
rect 15406 20194 15440 20228
rect 15406 20126 15440 20160
rect 15406 20058 15440 20092
rect 15406 19990 15440 20024
rect 15406 19922 15440 19956
rect 15406 19854 15440 19888
rect 15406 19786 15440 19820
rect 15406 19718 15440 19752
rect 15406 19650 15440 19684
rect 15406 19582 15440 19616
rect 15406 19514 15440 19548
rect 15406 19446 15440 19480
rect 15406 19378 15440 19412
rect 15406 19310 15440 19344
rect 15406 19242 15440 19276
rect 15406 19174 15440 19208
rect 15502 20398 15536 20432
rect 15502 20330 15536 20364
rect 15502 20262 15536 20296
rect 15502 20194 15536 20228
rect 15502 20126 15536 20160
rect 15502 20058 15536 20092
rect 15502 19990 15536 20024
rect 15502 19922 15536 19956
rect 15502 19854 15536 19888
rect 15502 19786 15536 19820
rect 15502 19718 15536 19752
rect 15502 19650 15536 19684
rect 15502 19582 15536 19616
rect 15502 19514 15536 19548
rect 15502 19446 15536 19480
rect 15502 19378 15536 19412
rect 15502 19310 15536 19344
rect 15502 19242 15536 19276
rect 15502 19174 15536 19208
rect 15990 19883 16024 19917
rect 15990 19815 16024 19849
rect 15990 19747 16024 19781
rect 15990 19679 16024 19713
rect 15990 19611 16024 19645
rect 15990 19543 16024 19577
rect 15990 19475 16024 19509
rect 15990 19407 16024 19441
rect 15990 19339 16024 19373
rect 15990 19271 16024 19305
rect 15990 19203 16024 19237
rect 16086 19883 16120 19917
rect 16086 19815 16120 19849
rect 16086 19747 16120 19781
rect 16086 19679 16120 19713
rect 16086 19611 16120 19645
rect 16086 19543 16120 19577
rect 16086 19475 16120 19509
rect 16086 19407 16120 19441
rect 16086 19339 16120 19373
rect 16086 19271 16120 19305
rect 16086 19203 16120 19237
rect 16182 19883 16216 19917
rect 16182 19815 16216 19849
rect 16182 19747 16216 19781
rect 16182 19679 16216 19713
rect 16182 19611 16216 19645
rect 16182 19543 16216 19577
rect 16182 19475 16216 19509
rect 16182 19407 16216 19441
rect 16182 19339 16216 19373
rect 16182 19271 16216 19305
rect 16182 19203 16216 19237
rect 16278 19883 16312 19917
rect 16278 19815 16312 19849
rect 16278 19747 16312 19781
rect 16278 19679 16312 19713
rect 16278 19611 16312 19645
rect 16278 19543 16312 19577
rect 16278 19475 16312 19509
rect 16278 19407 16312 19441
rect 16278 19339 16312 19373
rect 16278 19271 16312 19305
rect 16278 19203 16312 19237
rect 15016 18445 15050 18479
rect 15016 18377 15050 18411
rect 15016 18309 15050 18343
rect 15016 18241 15050 18275
rect 15016 18173 15050 18207
rect 15016 18105 15050 18139
rect 15016 18037 15050 18071
rect 15016 17969 15050 18003
rect 15016 17901 15050 17935
rect 15016 17833 15050 17867
rect 15016 17765 15050 17799
rect 15016 17697 15050 17731
rect 15016 17629 15050 17663
rect 15016 17561 15050 17595
rect 15016 17493 15050 17527
rect 15016 17425 15050 17459
rect 15016 17357 15050 17391
rect 15016 17289 15050 17323
rect 15016 17221 15050 17255
rect 15016 17153 15050 17187
rect 15016 17085 15050 17119
rect 15016 17017 15050 17051
rect 15016 16949 15050 16983
rect 15104 18445 15138 18479
rect 15104 18377 15138 18411
rect 15104 18309 15138 18343
rect 15104 18241 15138 18275
rect 15104 18173 15138 18207
rect 15104 18105 15138 18139
rect 15104 18037 15138 18071
rect 15104 17969 15138 18003
rect 15104 17901 15138 17935
rect 15104 17833 15138 17867
rect 15104 17765 15138 17799
rect 15104 17697 15138 17731
rect 15104 17629 15138 17663
rect 15104 17561 15138 17595
rect 15104 17493 15138 17527
rect 15104 17425 15138 17459
rect 15104 17357 15138 17391
rect 15104 17289 15138 17323
rect 15104 17221 15138 17255
rect 15104 17153 15138 17187
rect 15104 17085 15138 17119
rect 15104 17017 15138 17051
rect 15104 16949 15138 16983
rect 15426 18445 15460 18479
rect 15426 18377 15460 18411
rect 15426 18309 15460 18343
rect 15426 18241 15460 18275
rect 15426 18173 15460 18207
rect 15426 18105 15460 18139
rect 15426 18037 15460 18071
rect 15426 17969 15460 18003
rect 15426 17901 15460 17935
rect 15426 17833 15460 17867
rect 15426 17765 15460 17799
rect 15426 17697 15460 17731
rect 15426 17629 15460 17663
rect 15426 17561 15460 17595
rect 15426 17493 15460 17527
rect 15426 17425 15460 17459
rect 15426 17357 15460 17391
rect 15426 17289 15460 17323
rect 15426 17221 15460 17255
rect 15426 17153 15460 17187
rect 15426 17085 15460 17119
rect 15426 17017 15460 17051
rect 15426 16949 15460 16983
rect 15514 18445 15548 18479
rect 15514 18377 15548 18411
rect 15514 18309 15548 18343
rect 15514 18241 15548 18275
rect 15514 18173 15548 18207
rect 15514 18105 15548 18139
rect 15514 18037 15548 18071
rect 15514 17969 15548 18003
rect 15514 17901 15548 17935
rect 15514 17833 15548 17867
rect 15514 17765 15548 17799
rect 15514 17697 15548 17731
rect 15514 17629 15548 17663
rect 15514 17561 15548 17595
rect 15514 17493 15548 17527
rect 15514 17425 15548 17459
rect 15514 17357 15548 17391
rect 15514 17289 15548 17323
rect 15514 17221 15548 17255
rect 15514 17153 15548 17187
rect 15514 17085 15548 17119
rect 15514 17017 15548 17051
rect 15514 16949 15548 16983
rect 13572 15415 13606 15449
rect 13572 15347 13606 15381
rect 13572 15279 13606 15313
rect 13572 15211 13606 15245
rect 13572 15143 13606 15177
rect 13572 15075 13606 15109
rect 13572 15007 13606 15041
rect 13572 14939 13606 14973
rect 13572 14871 13606 14905
rect 13572 14803 13606 14837
rect 13572 14735 13606 14769
rect 13572 14667 13606 14701
rect 13572 14599 13606 14633
rect 13572 14531 13606 14565
rect 13572 14463 13606 14497
rect 13572 14395 13606 14429
rect 13572 14327 13606 14361
rect 13572 14259 13606 14293
rect 13572 14191 13606 14225
rect 13572 14123 13606 14157
rect 13572 14055 13606 14089
rect 13572 13987 13606 14021
rect 13572 13919 13606 13953
rect 13660 15415 13694 15449
rect 13660 15347 13694 15381
rect 13660 15279 13694 15313
rect 13660 15211 13694 15245
rect 13660 15143 13694 15177
rect 13660 15075 13694 15109
rect 13660 15007 13694 15041
rect 13660 14939 13694 14973
rect 13660 14871 13694 14905
rect 13660 14803 13694 14837
rect 13660 14735 13694 14769
rect 13660 14667 13694 14701
rect 13660 14599 13694 14633
rect 13660 14531 13694 14565
rect 13660 14463 13694 14497
rect 13660 14395 13694 14429
rect 13660 14327 13694 14361
rect 13660 14259 13694 14293
rect 13660 14191 13694 14225
rect 13660 14123 13694 14157
rect 13660 14055 13694 14089
rect 13660 13987 13694 14021
rect 13660 13919 13694 13953
rect 14422 15839 14456 15873
rect 14422 15771 14456 15805
rect 14422 15703 14456 15737
rect 14422 15635 14456 15669
rect 14422 15567 14456 15601
rect 14422 15499 14456 15533
rect 14422 15431 14456 15465
rect 14422 15363 14456 15397
rect 14422 15295 14456 15329
rect 14422 15227 14456 15261
rect 14422 15159 14456 15193
rect 14422 15091 14456 15125
rect 14422 15023 14456 15057
rect 14422 14955 14456 14989
rect 14422 14887 14456 14921
rect 14422 14819 14456 14853
rect 14422 14751 14456 14785
rect 14422 14683 14456 14717
rect 14422 14615 14456 14649
rect 14422 14547 14456 14581
rect 14422 14479 14456 14513
rect 14422 14411 14456 14445
rect 14422 14343 14456 14377
rect 14422 14275 14456 14309
rect 14422 14207 14456 14241
rect 14422 14139 14456 14173
rect 14422 14071 14456 14105
rect 14422 14003 14456 14037
rect 14422 13935 14456 13969
rect 14518 15839 14552 15873
rect 14518 15771 14552 15805
rect 14518 15703 14552 15737
rect 14518 15635 14552 15669
rect 14518 15567 14552 15601
rect 14518 15499 14552 15533
rect 14518 15431 14552 15465
rect 14518 15363 14552 15397
rect 14518 15295 14552 15329
rect 14518 15227 14552 15261
rect 14518 15159 14552 15193
rect 14518 15091 14552 15125
rect 14518 15023 14552 15057
rect 14518 14955 14552 14989
rect 14518 14887 14552 14921
rect 14518 14819 14552 14853
rect 14518 14751 14552 14785
rect 14518 14683 14552 14717
rect 14518 14615 14552 14649
rect 14518 14547 14552 14581
rect 14518 14479 14552 14513
rect 14518 14411 14552 14445
rect 14518 14343 14552 14377
rect 14518 14275 14552 14309
rect 14518 14207 14552 14241
rect 14518 14139 14552 14173
rect 14518 14071 14552 14105
rect 14518 14003 14552 14037
rect 14518 13935 14552 13969
rect 14614 15839 14648 15873
rect 14614 15771 14648 15805
rect 14614 15703 14648 15737
rect 14614 15635 14648 15669
rect 14614 15567 14648 15601
rect 14614 15499 14648 15533
rect 14614 15431 14648 15465
rect 14614 15363 14648 15397
rect 14614 15295 14648 15329
rect 14614 15227 14648 15261
rect 14614 15159 14648 15193
rect 14614 15091 14648 15125
rect 14614 15023 14648 15057
rect 14614 14955 14648 14989
rect 14614 14887 14648 14921
rect 14614 14819 14648 14853
rect 14614 14751 14648 14785
rect 14614 14683 14648 14717
rect 14614 14615 14648 14649
rect 14614 14547 14648 14581
rect 14614 14479 14648 14513
rect 14614 14411 14648 14445
rect 14614 14343 14648 14377
rect 14614 14275 14648 14309
rect 14614 14207 14648 14241
rect 14614 14139 14648 14173
rect 14614 14071 14648 14105
rect 14614 14003 14648 14037
rect 14614 13935 14648 13969
rect 14710 15839 14744 15873
rect 14710 15771 14744 15805
rect 14710 15703 14744 15737
rect 14710 15635 14744 15669
rect 14710 15567 14744 15601
rect 14710 15499 14744 15533
rect 14710 15431 14744 15465
rect 14710 15363 14744 15397
rect 14710 15295 14744 15329
rect 14710 15227 14744 15261
rect 14710 15159 14744 15193
rect 14710 15091 14744 15125
rect 14710 15023 14744 15057
rect 14710 14955 14744 14989
rect 14710 14887 14744 14921
rect 14710 14819 14744 14853
rect 14710 14751 14744 14785
rect 14710 14683 14744 14717
rect 14710 14615 14744 14649
rect 14710 14547 14744 14581
rect 14710 14479 14744 14513
rect 14710 14411 14744 14445
rect 14710 14343 14744 14377
rect 14710 14275 14744 14309
rect 14710 14207 14744 14241
rect 14710 14139 14744 14173
rect 14710 14071 14744 14105
rect 14710 14003 14744 14037
rect 14710 13935 14744 13969
rect 14806 15839 14840 15873
rect 14806 15771 14840 15805
rect 14806 15703 14840 15737
rect 14806 15635 14840 15669
rect 14806 15567 14840 15601
rect 14806 15499 14840 15533
rect 14806 15431 14840 15465
rect 14806 15363 14840 15397
rect 14806 15295 14840 15329
rect 14806 15227 14840 15261
rect 14806 15159 14840 15193
rect 14806 15091 14840 15125
rect 14806 15023 14840 15057
rect 14806 14955 14840 14989
rect 14806 14887 14840 14921
rect 14806 14819 14840 14853
rect 14806 14751 14840 14785
rect 14806 14683 14840 14717
rect 14806 14615 14840 14649
rect 14806 14547 14840 14581
rect 14806 14479 14840 14513
rect 14806 14411 14840 14445
rect 14806 14343 14840 14377
rect 14806 14275 14840 14309
rect 14806 14207 14840 14241
rect 14806 14139 14840 14173
rect 14806 14071 14840 14105
rect 14806 14003 14840 14037
rect 14806 13935 14840 13969
rect 14902 15839 14936 15873
rect 14902 15771 14936 15805
rect 14902 15703 14936 15737
rect 14902 15635 14936 15669
rect 14902 15567 14936 15601
rect 14902 15499 14936 15533
rect 14902 15431 14936 15465
rect 14902 15363 14936 15397
rect 14902 15295 14936 15329
rect 14902 15227 14936 15261
rect 14902 15159 14936 15193
rect 14902 15091 14936 15125
rect 14902 15023 14936 15057
rect 14902 14955 14936 14989
rect 14902 14887 14936 14921
rect 14902 14819 14936 14853
rect 14902 14751 14936 14785
rect 14902 14683 14936 14717
rect 14902 14615 14936 14649
rect 14902 14547 14936 14581
rect 14902 14479 14936 14513
rect 14902 14411 14936 14445
rect 14902 14343 14936 14377
rect 14902 14275 14936 14309
rect 14902 14207 14936 14241
rect 14902 14139 14936 14173
rect 14902 14071 14936 14105
rect 14902 14003 14936 14037
rect 14902 13935 14936 13969
rect 14998 15839 15032 15873
rect 14998 15771 15032 15805
rect 14998 15703 15032 15737
rect 14998 15635 15032 15669
rect 14998 15567 15032 15601
rect 14998 15499 15032 15533
rect 14998 15431 15032 15465
rect 14998 15363 15032 15397
rect 14998 15295 15032 15329
rect 14998 15227 15032 15261
rect 14998 15159 15032 15193
rect 14998 15091 15032 15125
rect 14998 15023 15032 15057
rect 14998 14955 15032 14989
rect 14998 14887 15032 14921
rect 14998 14819 15032 14853
rect 14998 14751 15032 14785
rect 14998 14683 15032 14717
rect 14998 14615 15032 14649
rect 14998 14547 15032 14581
rect 14998 14479 15032 14513
rect 14998 14411 15032 14445
rect 14998 14343 15032 14377
rect 14998 14275 15032 14309
rect 14998 14207 15032 14241
rect 14998 14139 15032 14173
rect 14998 14071 15032 14105
rect 14998 14003 15032 14037
rect 14998 13935 15032 13969
rect 15094 15839 15128 15873
rect 15094 15771 15128 15805
rect 15094 15703 15128 15737
rect 15094 15635 15128 15669
rect 15094 15567 15128 15601
rect 15094 15499 15128 15533
rect 15094 15431 15128 15465
rect 15094 15363 15128 15397
rect 15094 15295 15128 15329
rect 15094 15227 15128 15261
rect 15094 15159 15128 15193
rect 15094 15091 15128 15125
rect 15094 15023 15128 15057
rect 15094 14955 15128 14989
rect 15094 14887 15128 14921
rect 15094 14819 15128 14853
rect 15094 14751 15128 14785
rect 15094 14683 15128 14717
rect 15094 14615 15128 14649
rect 15094 14547 15128 14581
rect 15094 14479 15128 14513
rect 15094 14411 15128 14445
rect 15094 14343 15128 14377
rect 15094 14275 15128 14309
rect 15094 14207 15128 14241
rect 15094 14139 15128 14173
rect 15094 14071 15128 14105
rect 15094 14003 15128 14037
rect 15094 13935 15128 13969
rect 15190 15839 15224 15873
rect 15190 15771 15224 15805
rect 15190 15703 15224 15737
rect 15190 15635 15224 15669
rect 15190 15567 15224 15601
rect 15190 15499 15224 15533
rect 15190 15431 15224 15465
rect 15190 15363 15224 15397
rect 15190 15295 15224 15329
rect 15190 15227 15224 15261
rect 15190 15159 15224 15193
rect 15190 15091 15224 15125
rect 15190 15023 15224 15057
rect 15190 14955 15224 14989
rect 15190 14887 15224 14921
rect 15190 14819 15224 14853
rect 15190 14751 15224 14785
rect 15190 14683 15224 14717
rect 15190 14615 15224 14649
rect 15190 14547 15224 14581
rect 15190 14479 15224 14513
rect 15190 14411 15224 14445
rect 15190 14343 15224 14377
rect 15190 14275 15224 14309
rect 15190 14207 15224 14241
rect 15190 14139 15224 14173
rect 15190 14071 15224 14105
rect 15190 14003 15224 14037
rect 15190 13935 15224 13969
rect 13434 13005 13468 13039
rect 13434 12937 13468 12971
rect 13434 12869 13468 12903
rect 13434 12801 13468 12835
rect 13434 12733 13468 12767
rect 13434 12665 13468 12699
rect 13434 12597 13468 12631
rect 13434 12529 13468 12563
rect 13434 12461 13468 12495
rect 13434 12393 13468 12427
rect 13434 12325 13468 12359
rect 13434 12257 13468 12291
rect 13434 12189 13468 12223
rect 13434 12121 13468 12155
rect 13434 12053 13468 12087
rect 13434 11985 13468 12019
rect 13434 11917 13468 11951
rect 13434 11849 13468 11883
rect 13434 11781 13468 11815
rect 13434 11713 13468 11747
rect 13434 11645 13468 11679
rect 13434 11577 13468 11611
rect 13434 11509 13468 11543
rect 13434 11441 13468 11475
rect 13434 11373 13468 11407
rect 13434 11305 13468 11339
rect 13434 11237 13468 11271
rect 13434 11169 13468 11203
rect 13434 11101 13468 11135
rect 13522 13005 13556 13039
rect 13522 12937 13556 12971
rect 13522 12869 13556 12903
rect 13522 12801 13556 12835
rect 13522 12733 13556 12767
rect 13522 12665 13556 12699
rect 13522 12597 13556 12631
rect 13522 12529 13556 12563
rect 13522 12461 13556 12495
rect 13522 12393 13556 12427
rect 13522 12325 13556 12359
rect 13522 12257 13556 12291
rect 13522 12189 13556 12223
rect 13522 12121 13556 12155
rect 13522 12053 13556 12087
rect 13522 11985 13556 12019
rect 13522 11917 13556 11951
rect 13522 11849 13556 11883
rect 13522 11781 13556 11815
rect 13522 11713 13556 11747
rect 13522 11645 13556 11679
rect 13522 11577 13556 11611
rect 13522 11509 13556 11543
rect 13522 11441 13556 11475
rect 13522 11373 13556 11407
rect 13522 11305 13556 11339
rect 13522 11237 13556 11271
rect 13522 11169 13556 11203
rect 13522 11101 13556 11135
rect 13610 13005 13644 13039
rect 13610 12937 13644 12971
rect 13610 12869 13644 12903
rect 13610 12801 13644 12835
rect 13610 12733 13644 12767
rect 13610 12665 13644 12699
rect 13610 12597 13644 12631
rect 13610 12529 13644 12563
rect 13610 12461 13644 12495
rect 13610 12393 13644 12427
rect 13610 12325 13644 12359
rect 13610 12257 13644 12291
rect 13610 12189 13644 12223
rect 13610 12121 13644 12155
rect 13610 12053 13644 12087
rect 13610 11985 13644 12019
rect 13610 11917 13644 11951
rect 13610 11849 13644 11883
rect 13610 11781 13644 11815
rect 13610 11713 13644 11747
rect 13610 11645 13644 11679
rect 13610 11577 13644 11611
rect 13610 11509 13644 11543
rect 13610 11441 13644 11475
rect 13610 11373 13644 11407
rect 13610 11305 13644 11339
rect 13610 11237 13644 11271
rect 13610 11169 13644 11203
rect 13610 11101 13644 11135
rect 13698 13005 13732 13039
rect 13698 12937 13732 12971
rect 13698 12869 13732 12903
rect 13698 12801 13732 12835
rect 13698 12733 13732 12767
rect 13698 12665 13732 12699
rect 13698 12597 13732 12631
rect 13698 12529 13732 12563
rect 13698 12461 13732 12495
rect 13698 12393 13732 12427
rect 13698 12325 13732 12359
rect 13698 12257 13732 12291
rect 13698 12189 13732 12223
rect 13698 12121 13732 12155
rect 13698 12053 13732 12087
rect 13698 11985 13732 12019
rect 13698 11917 13732 11951
rect 13698 11849 13732 11883
rect 13698 11781 13732 11815
rect 13698 11713 13732 11747
rect 13698 11645 13732 11679
rect 13698 11577 13732 11611
rect 13698 11509 13732 11543
rect 13698 11441 13732 11475
rect 13698 11373 13732 11407
rect 13698 11305 13732 11339
rect 13698 11237 13732 11271
rect 13698 11169 13732 11203
rect 13698 11101 13732 11135
rect 13786 13005 13820 13039
rect 13786 12937 13820 12971
rect 13786 12869 13820 12903
rect 13786 12801 13820 12835
rect 13786 12733 13820 12767
rect 13786 12665 13820 12699
rect 13786 12597 13820 12631
rect 13786 12529 13820 12563
rect 13786 12461 13820 12495
rect 13786 12393 13820 12427
rect 13786 12325 13820 12359
rect 13786 12257 13820 12291
rect 13786 12189 13820 12223
rect 13786 12121 13820 12155
rect 13786 12053 13820 12087
rect 13786 11985 13820 12019
rect 13786 11917 13820 11951
rect 13786 11849 13820 11883
rect 13786 11781 13820 11815
rect 13786 11713 13820 11747
rect 13786 11645 13820 11679
rect 13786 11577 13820 11611
rect 13786 11509 13820 11543
rect 13786 11441 13820 11475
rect 13786 11373 13820 11407
rect 13786 11305 13820 11339
rect 13786 11237 13820 11271
rect 13786 11169 13820 11203
rect 13786 11101 13820 11135
rect 13874 13005 13908 13039
rect 13874 12937 13908 12971
rect 13874 12869 13908 12903
rect 13874 12801 13908 12835
rect 13874 12733 13908 12767
rect 13874 12665 13908 12699
rect 13874 12597 13908 12631
rect 13874 12529 13908 12563
rect 13874 12461 13908 12495
rect 13874 12393 13908 12427
rect 13874 12325 13908 12359
rect 13874 12257 13908 12291
rect 13874 12189 13908 12223
rect 13874 12121 13908 12155
rect 13874 12053 13908 12087
rect 13874 11985 13908 12019
rect 13874 11917 13908 11951
rect 13874 11849 13908 11883
rect 13874 11781 13908 11815
rect 13874 11713 13908 11747
rect 13874 11645 13908 11679
rect 13874 11577 13908 11611
rect 13874 11509 13908 11543
rect 13874 11441 13908 11475
rect 13874 11373 13908 11407
rect 13874 11305 13908 11339
rect 13874 11237 13908 11271
rect 13874 11169 13908 11203
rect 13874 11101 13908 11135
rect 13962 13005 13996 13039
rect 13962 12937 13996 12971
rect 13962 12869 13996 12903
rect 13962 12801 13996 12835
rect 13962 12733 13996 12767
rect 13962 12665 13996 12699
rect 13962 12597 13996 12631
rect 13962 12529 13996 12563
rect 13962 12461 13996 12495
rect 13962 12393 13996 12427
rect 13962 12325 13996 12359
rect 13962 12257 13996 12291
rect 13962 12189 13996 12223
rect 13962 12121 13996 12155
rect 13962 12053 13996 12087
rect 13962 11985 13996 12019
rect 13962 11917 13996 11951
rect 13962 11849 13996 11883
rect 13962 11781 13996 11815
rect 13962 11713 13996 11747
rect 13962 11645 13996 11679
rect 13962 11577 13996 11611
rect 13962 11509 13996 11543
rect 13962 11441 13996 11475
rect 13962 11373 13996 11407
rect 13962 11305 13996 11339
rect 13962 11237 13996 11271
rect 13962 11169 13996 11203
rect 13962 11101 13996 11135
rect 14050 13005 14084 13039
rect 14050 12937 14084 12971
rect 14050 12869 14084 12903
rect 14050 12801 14084 12835
rect 14050 12733 14084 12767
rect 14050 12665 14084 12699
rect 14050 12597 14084 12631
rect 14050 12529 14084 12563
rect 14050 12461 14084 12495
rect 14050 12393 14084 12427
rect 14050 12325 14084 12359
rect 14050 12257 14084 12291
rect 14050 12189 14084 12223
rect 14050 12121 14084 12155
rect 14050 12053 14084 12087
rect 14050 11985 14084 12019
rect 14050 11917 14084 11951
rect 14050 11849 14084 11883
rect 14050 11781 14084 11815
rect 14050 11713 14084 11747
rect 14050 11645 14084 11679
rect 14050 11577 14084 11611
rect 14050 11509 14084 11543
rect 14050 11441 14084 11475
rect 14050 11373 14084 11407
rect 14050 11305 14084 11339
rect 14050 11237 14084 11271
rect 14050 11169 14084 11203
rect 14050 11101 14084 11135
rect 14138 13005 14172 13039
rect 14138 12937 14172 12971
rect 14138 12869 14172 12903
rect 14138 12801 14172 12835
rect 14138 12733 14172 12767
rect 14138 12665 14172 12699
rect 14138 12597 14172 12631
rect 14138 12529 14172 12563
rect 14138 12461 14172 12495
rect 14138 12393 14172 12427
rect 14138 12325 14172 12359
rect 14138 12257 14172 12291
rect 14138 12189 14172 12223
rect 14138 12121 14172 12155
rect 14138 12053 14172 12087
rect 14138 11985 14172 12019
rect 14138 11917 14172 11951
rect 14138 11849 14172 11883
rect 14138 11781 14172 11815
rect 14138 11713 14172 11747
rect 14138 11645 14172 11679
rect 14138 11577 14172 11611
rect 14138 11509 14172 11543
rect 14138 11441 14172 11475
rect 14138 11373 14172 11407
rect 14138 11305 14172 11339
rect 14138 11237 14172 11271
rect 14138 11169 14172 11203
rect 14138 11101 14172 11135
rect 14226 13005 14260 13039
rect 14226 12937 14260 12971
rect 14226 12869 14260 12903
rect 14226 12801 14260 12835
rect 14226 12733 14260 12767
rect 14226 12665 14260 12699
rect 14226 12597 14260 12631
rect 14226 12529 14260 12563
rect 14226 12461 14260 12495
rect 14226 12393 14260 12427
rect 14226 12325 14260 12359
rect 14226 12257 14260 12291
rect 14226 12189 14260 12223
rect 14226 12121 14260 12155
rect 14226 12053 14260 12087
rect 14226 11985 14260 12019
rect 14226 11917 14260 11951
rect 14226 11849 14260 11883
rect 14226 11781 14260 11815
rect 14226 11713 14260 11747
rect 14226 11645 14260 11679
rect 14226 11577 14260 11611
rect 14226 11509 14260 11543
rect 14226 11441 14260 11475
rect 14226 11373 14260 11407
rect 14226 11305 14260 11339
rect 14226 11237 14260 11271
rect 14226 11169 14260 11203
rect 14226 11101 14260 11135
rect 14314 13005 14348 13039
rect 14314 12937 14348 12971
rect 14314 12869 14348 12903
rect 14314 12801 14348 12835
rect 14314 12733 14348 12767
rect 14314 12665 14348 12699
rect 14314 12597 14348 12631
rect 14314 12529 14348 12563
rect 14314 12461 14348 12495
rect 14314 12393 14348 12427
rect 14314 12325 14348 12359
rect 14314 12257 14348 12291
rect 14314 12189 14348 12223
rect 14314 12121 14348 12155
rect 14314 12053 14348 12087
rect 14314 11985 14348 12019
rect 14314 11917 14348 11951
rect 14314 11849 14348 11883
rect 14314 11781 14348 11815
rect 14314 11713 14348 11747
rect 14314 11645 14348 11679
rect 14314 11577 14348 11611
rect 14314 11509 14348 11543
rect 14314 11441 14348 11475
rect 14314 11373 14348 11407
rect 14314 11305 14348 11339
rect 14314 11237 14348 11271
rect 14314 11169 14348 11203
rect 14314 11101 14348 11135
rect 14402 13005 14436 13039
rect 14402 12937 14436 12971
rect 14402 12869 14436 12903
rect 14402 12801 14436 12835
rect 14402 12733 14436 12767
rect 14402 12665 14436 12699
rect 14402 12597 14436 12631
rect 14402 12529 14436 12563
rect 14402 12461 14436 12495
rect 14402 12393 14436 12427
rect 14402 12325 14436 12359
rect 14402 12257 14436 12291
rect 14402 12189 14436 12223
rect 14402 12121 14436 12155
rect 14402 12053 14436 12087
rect 14402 11985 14436 12019
rect 14402 11917 14436 11951
rect 14402 11849 14436 11883
rect 14402 11781 14436 11815
rect 14402 11713 14436 11747
rect 14402 11645 14436 11679
rect 14402 11577 14436 11611
rect 14402 11509 14436 11543
rect 14402 11441 14436 11475
rect 14402 11373 14436 11407
rect 14402 11305 14436 11339
rect 14402 11237 14436 11271
rect 14402 11169 14436 11203
rect 14402 11101 14436 11135
rect 14490 13005 14524 13039
rect 14490 12937 14524 12971
rect 14490 12869 14524 12903
rect 14490 12801 14524 12835
rect 14490 12733 14524 12767
rect 14490 12665 14524 12699
rect 14490 12597 14524 12631
rect 14490 12529 14524 12563
rect 14490 12461 14524 12495
rect 14490 12393 14524 12427
rect 14490 12325 14524 12359
rect 14490 12257 14524 12291
rect 14490 12189 14524 12223
rect 14490 12121 14524 12155
rect 14490 12053 14524 12087
rect 14490 11985 14524 12019
rect 14490 11917 14524 11951
rect 14490 11849 14524 11883
rect 14490 11781 14524 11815
rect 14490 11713 14524 11747
rect 14490 11645 14524 11679
rect 14490 11577 14524 11611
rect 14490 11509 14524 11543
rect 14490 11441 14524 11475
rect 14490 11373 14524 11407
rect 14490 11305 14524 11339
rect 14490 11237 14524 11271
rect 14490 11169 14524 11203
rect 14490 11101 14524 11135
rect 14578 13005 14612 13039
rect 14578 12937 14612 12971
rect 14578 12869 14612 12903
rect 14578 12801 14612 12835
rect 14578 12733 14612 12767
rect 14578 12665 14612 12699
rect 14578 12597 14612 12631
rect 14578 12529 14612 12563
rect 14578 12461 14612 12495
rect 14578 12393 14612 12427
rect 14578 12325 14612 12359
rect 14578 12257 14612 12291
rect 14578 12189 14612 12223
rect 14578 12121 14612 12155
rect 14578 12053 14612 12087
rect 14578 11985 14612 12019
rect 14578 11917 14612 11951
rect 14578 11849 14612 11883
rect 14578 11781 14612 11815
rect 14578 11713 14612 11747
rect 14578 11645 14612 11679
rect 14578 11577 14612 11611
rect 14578 11509 14612 11543
rect 14578 11441 14612 11475
rect 14578 11373 14612 11407
rect 14578 11305 14612 11339
rect 14578 11237 14612 11271
rect 14578 11169 14612 11203
rect 14578 11101 14612 11135
rect 14666 13005 14700 13039
rect 14666 12937 14700 12971
rect 14666 12869 14700 12903
rect 14666 12801 14700 12835
rect 14666 12733 14700 12767
rect 14666 12665 14700 12699
rect 14666 12597 14700 12631
rect 14666 12529 14700 12563
rect 14666 12461 14700 12495
rect 14666 12393 14700 12427
rect 14666 12325 14700 12359
rect 14666 12257 14700 12291
rect 14666 12189 14700 12223
rect 14666 12121 14700 12155
rect 14666 12053 14700 12087
rect 14666 11985 14700 12019
rect 14666 11917 14700 11951
rect 14666 11849 14700 11883
rect 14666 11781 14700 11815
rect 14666 11713 14700 11747
rect 14666 11645 14700 11679
rect 14666 11577 14700 11611
rect 14666 11509 14700 11543
rect 14666 11441 14700 11475
rect 14666 11373 14700 11407
rect 14666 11305 14700 11339
rect 14666 11237 14700 11271
rect 14666 11169 14700 11203
rect 14666 11101 14700 11135
rect 14754 13005 14788 13039
rect 14754 12937 14788 12971
rect 14754 12869 14788 12903
rect 14754 12801 14788 12835
rect 14754 12733 14788 12767
rect 14754 12665 14788 12699
rect 14754 12597 14788 12631
rect 14754 12529 14788 12563
rect 14754 12461 14788 12495
rect 14754 12393 14788 12427
rect 14754 12325 14788 12359
rect 14754 12257 14788 12291
rect 14754 12189 14788 12223
rect 14754 12121 14788 12155
rect 14754 12053 14788 12087
rect 14754 11985 14788 12019
rect 14754 11917 14788 11951
rect 14754 11849 14788 11883
rect 14754 11781 14788 11815
rect 14754 11713 14788 11747
rect 14754 11645 14788 11679
rect 14754 11577 14788 11611
rect 14754 11509 14788 11543
rect 14754 11441 14788 11475
rect 14754 11373 14788 11407
rect 14754 11305 14788 11339
rect 14754 11237 14788 11271
rect 14754 11169 14788 11203
rect 14754 11101 14788 11135
rect 14842 13005 14876 13039
rect 14842 12937 14876 12971
rect 14842 12869 14876 12903
rect 14842 12801 14876 12835
rect 14842 12733 14876 12767
rect 14842 12665 14876 12699
rect 14842 12597 14876 12631
rect 14842 12529 14876 12563
rect 14842 12461 14876 12495
rect 14842 12393 14876 12427
rect 14842 12325 14876 12359
rect 14842 12257 14876 12291
rect 14842 12189 14876 12223
rect 14842 12121 14876 12155
rect 14842 12053 14876 12087
rect 14842 11985 14876 12019
rect 14842 11917 14876 11951
rect 14842 11849 14876 11883
rect 14842 11781 14876 11815
rect 14842 11713 14876 11747
rect 14842 11645 14876 11679
rect 14842 11577 14876 11611
rect 14842 11509 14876 11543
rect 14842 11441 14876 11475
rect 14842 11373 14876 11407
rect 14842 11305 14876 11339
rect 14842 11237 14876 11271
rect 14842 11169 14876 11203
rect 14842 11101 14876 11135
rect 14930 13005 14964 13039
rect 14930 12937 14964 12971
rect 14930 12869 14964 12903
rect 14930 12801 14964 12835
rect 14930 12733 14964 12767
rect 14930 12665 14964 12699
rect 14930 12597 14964 12631
rect 14930 12529 14964 12563
rect 14930 12461 14964 12495
rect 14930 12393 14964 12427
rect 14930 12325 14964 12359
rect 14930 12257 14964 12291
rect 14930 12189 14964 12223
rect 14930 12121 14964 12155
rect 14930 12053 14964 12087
rect 14930 11985 14964 12019
rect 14930 11917 14964 11951
rect 14930 11849 14964 11883
rect 14930 11781 14964 11815
rect 14930 11713 14964 11747
rect 14930 11645 14964 11679
rect 14930 11577 14964 11611
rect 14930 11509 14964 11543
rect 14930 11441 14964 11475
rect 14930 11373 14964 11407
rect 14930 11305 14964 11339
rect 14930 11237 14964 11271
rect 14930 11169 14964 11203
rect 14930 11101 14964 11135
rect 15018 13005 15052 13039
rect 15018 12937 15052 12971
rect 15018 12869 15052 12903
rect 15018 12801 15052 12835
rect 15018 12733 15052 12767
rect 15018 12665 15052 12699
rect 15018 12597 15052 12631
rect 15018 12529 15052 12563
rect 15018 12461 15052 12495
rect 15018 12393 15052 12427
rect 15018 12325 15052 12359
rect 15018 12257 15052 12291
rect 15018 12189 15052 12223
rect 15018 12121 15052 12155
rect 15018 12053 15052 12087
rect 15018 11985 15052 12019
rect 15018 11917 15052 11951
rect 15018 11849 15052 11883
rect 15018 11781 15052 11815
rect 15018 11713 15052 11747
rect 15018 11645 15052 11679
rect 15018 11577 15052 11611
rect 15018 11509 15052 11543
rect 15018 11441 15052 11475
rect 15018 11373 15052 11407
rect 15018 11305 15052 11339
rect 15018 11237 15052 11271
rect 15018 11169 15052 11203
rect 15018 11101 15052 11135
rect 15106 13005 15140 13039
rect 15106 12937 15140 12971
rect 15106 12869 15140 12903
rect 15106 12801 15140 12835
rect 15106 12733 15140 12767
rect 15106 12665 15140 12699
rect 15106 12597 15140 12631
rect 15106 12529 15140 12563
rect 15106 12461 15140 12495
rect 15106 12393 15140 12427
rect 15106 12325 15140 12359
rect 15106 12257 15140 12291
rect 15106 12189 15140 12223
rect 15106 12121 15140 12155
rect 15106 12053 15140 12087
rect 15106 11985 15140 12019
rect 15106 11917 15140 11951
rect 15106 11849 15140 11883
rect 15106 11781 15140 11815
rect 15106 11713 15140 11747
rect 15106 11645 15140 11679
rect 15106 11577 15140 11611
rect 15106 11509 15140 11543
rect 15106 11441 15140 11475
rect 15106 11373 15140 11407
rect 15106 11305 15140 11339
rect 15106 11237 15140 11271
rect 15106 11169 15140 11203
rect 15106 11101 15140 11135
rect 15194 13005 15228 13039
rect 15194 12937 15228 12971
rect 15194 12869 15228 12903
rect 15194 12801 15228 12835
rect 15194 12733 15228 12767
rect 15194 12665 15228 12699
rect 15194 12597 15228 12631
rect 15194 12529 15228 12563
rect 15194 12461 15228 12495
rect 15194 12393 15228 12427
rect 15194 12325 15228 12359
rect 15194 12257 15228 12291
rect 15194 12189 15228 12223
rect 15194 12121 15228 12155
rect 15194 12053 15228 12087
rect 15194 11985 15228 12019
rect 15194 11917 15228 11951
rect 15194 11849 15228 11883
rect 15194 11781 15228 11815
rect 15194 11713 15228 11747
rect 15194 11645 15228 11679
rect 15194 11577 15228 11611
rect 15194 11509 15228 11543
rect 15194 11441 15228 11475
rect 15194 11373 15228 11407
rect 15194 11305 15228 11339
rect 15194 11237 15228 11271
rect 15194 11169 15228 11203
rect 15194 11101 15228 11135
rect 15282 13005 15316 13039
rect 15282 12937 15316 12971
rect 15282 12869 15316 12903
rect 15282 12801 15316 12835
rect 15282 12733 15316 12767
rect 15282 12665 15316 12699
rect 15282 12597 15316 12631
rect 15282 12529 15316 12563
rect 15282 12461 15316 12495
rect 15282 12393 15316 12427
rect 15282 12325 15316 12359
rect 15282 12257 15316 12291
rect 15282 12189 15316 12223
rect 15282 12121 15316 12155
rect 15282 12053 15316 12087
rect 15282 11985 15316 12019
rect 15282 11917 15316 11951
rect 15282 11849 15316 11883
rect 15282 11781 15316 11815
rect 15282 11713 15316 11747
rect 15282 11645 15316 11679
rect 15282 11577 15316 11611
rect 15282 11509 15316 11543
rect 15282 11441 15316 11475
rect 15282 11373 15316 11407
rect 15282 11305 15316 11339
rect 15282 11237 15316 11271
rect 15282 11169 15316 11203
rect 15282 11101 15316 11135
rect 15370 13005 15404 13039
rect 15370 12937 15404 12971
rect 15370 12869 15404 12903
rect 15370 12801 15404 12835
rect 15370 12733 15404 12767
rect 15370 12665 15404 12699
rect 15370 12597 15404 12631
rect 15370 12529 15404 12563
rect 15370 12461 15404 12495
rect 15370 12393 15404 12427
rect 15370 12325 15404 12359
rect 15370 12257 15404 12291
rect 15370 12189 15404 12223
rect 15370 12121 15404 12155
rect 15370 12053 15404 12087
rect 15370 11985 15404 12019
rect 15370 11917 15404 11951
rect 15370 11849 15404 11883
rect 15370 11781 15404 11815
rect 15370 11713 15404 11747
rect 15370 11645 15404 11679
rect 15370 11577 15404 11611
rect 15370 11509 15404 11543
rect 15370 11441 15404 11475
rect 15370 11373 15404 11407
rect 15370 11305 15404 11339
rect 15370 11237 15404 11271
rect 15370 11169 15404 11203
rect 15370 11101 15404 11135
rect 15458 13005 15492 13039
rect 15458 12937 15492 12971
rect 15458 12869 15492 12903
rect 15458 12801 15492 12835
rect 15458 12733 15492 12767
rect 15458 12665 15492 12699
rect 15458 12597 15492 12631
rect 15458 12529 15492 12563
rect 15458 12461 15492 12495
rect 15458 12393 15492 12427
rect 15458 12325 15492 12359
rect 15458 12257 15492 12291
rect 15458 12189 15492 12223
rect 15458 12121 15492 12155
rect 15458 12053 15492 12087
rect 15458 11985 15492 12019
rect 15458 11917 15492 11951
rect 15458 11849 15492 11883
rect 15458 11781 15492 11815
rect 15458 11713 15492 11747
rect 15458 11645 15492 11679
rect 15458 11577 15492 11611
rect 15458 11509 15492 11543
rect 15458 11441 15492 11475
rect 15458 11373 15492 11407
rect 15458 11305 15492 11339
rect 15458 11237 15492 11271
rect 15458 11169 15492 11203
rect 15458 11101 15492 11135
rect 15546 13005 15580 13039
rect 15546 12937 15580 12971
rect 15546 12869 15580 12903
rect 15546 12801 15580 12835
rect 15546 12733 15580 12767
rect 15546 12665 15580 12699
rect 15546 12597 15580 12631
rect 15546 12529 15580 12563
rect 15546 12461 15580 12495
rect 15546 12393 15580 12427
rect 15546 12325 15580 12359
rect 15546 12257 15580 12291
rect 15546 12189 15580 12223
rect 15546 12121 15580 12155
rect 15546 12053 15580 12087
rect 15546 11985 15580 12019
rect 15546 11917 15580 11951
rect 15546 11849 15580 11883
rect 15546 11781 15580 11815
rect 15546 11713 15580 11747
rect 15546 11645 15580 11679
rect 15546 11577 15580 11611
rect 15546 11509 15580 11543
rect 15546 11441 15580 11475
rect 15546 11373 15580 11407
rect 15546 11305 15580 11339
rect 15546 11237 15580 11271
rect 15546 11169 15580 11203
rect 15546 11101 15580 11135
rect 15634 13005 15668 13039
rect 15634 12937 15668 12971
rect 15634 12869 15668 12903
rect 15634 12801 15668 12835
rect 15634 12733 15668 12767
rect 15634 12665 15668 12699
rect 15634 12597 15668 12631
rect 15634 12529 15668 12563
rect 15634 12461 15668 12495
rect 15634 12393 15668 12427
rect 15634 12325 15668 12359
rect 15634 12257 15668 12291
rect 15634 12189 15668 12223
rect 15634 12121 15668 12155
rect 15634 12053 15668 12087
rect 15634 11985 15668 12019
rect 15634 11917 15668 11951
rect 15634 11849 15668 11883
rect 15634 11781 15668 11815
rect 15634 11713 15668 11747
rect 15634 11645 15668 11679
rect 15634 11577 15668 11611
rect 15634 11509 15668 11543
rect 15634 11441 15668 11475
rect 15634 11373 15668 11407
rect 15634 11305 15668 11339
rect 15634 11237 15668 11271
rect 15634 11169 15668 11203
rect 15634 11101 15668 11135
rect 15722 13005 15756 13039
rect 15722 12937 15756 12971
rect 15722 12869 15756 12903
rect 15722 12801 15756 12835
rect 15722 12733 15756 12767
rect 15722 12665 15756 12699
rect 15722 12597 15756 12631
rect 15722 12529 15756 12563
rect 15722 12461 15756 12495
rect 15722 12393 15756 12427
rect 15722 12325 15756 12359
rect 15722 12257 15756 12291
rect 15722 12189 15756 12223
rect 15722 12121 15756 12155
rect 15722 12053 15756 12087
rect 15722 11985 15756 12019
rect 15722 11917 15756 11951
rect 15722 11849 15756 11883
rect 15722 11781 15756 11815
rect 15722 11713 15756 11747
rect 15722 11645 15756 11679
rect 15722 11577 15756 11611
rect 15722 11509 15756 11543
rect 15722 11441 15756 11475
rect 15722 11373 15756 11407
rect 15722 11305 15756 11339
rect 15722 11237 15756 11271
rect 15722 11169 15756 11203
rect 15722 11101 15756 11135
rect 15810 13005 15844 13039
rect 15810 12937 15844 12971
rect 15810 12869 15844 12903
rect 15810 12801 15844 12835
rect 15810 12733 15844 12767
rect 15810 12665 15844 12699
rect 15810 12597 15844 12631
rect 15810 12529 15844 12563
rect 15810 12461 15844 12495
rect 15810 12393 15844 12427
rect 15810 12325 15844 12359
rect 15810 12257 15844 12291
rect 15810 12189 15844 12223
rect 15810 12121 15844 12155
rect 15810 12053 15844 12087
rect 15810 11985 15844 12019
rect 15810 11917 15844 11951
rect 15810 11849 15844 11883
rect 15810 11781 15844 11815
rect 15810 11713 15844 11747
rect 15810 11645 15844 11679
rect 15810 11577 15844 11611
rect 15810 11509 15844 11543
rect 15810 11441 15844 11475
rect 15810 11373 15844 11407
rect 15810 11305 15844 11339
rect 15810 11237 15844 11271
rect 15810 11169 15844 11203
rect 15810 11101 15844 11135
rect 15898 13005 15932 13039
rect 15898 12937 15932 12971
rect 15898 12869 15932 12903
rect 15898 12801 15932 12835
rect 15898 12733 15932 12767
rect 15898 12665 15932 12699
rect 15898 12597 15932 12631
rect 15898 12529 15932 12563
rect 15898 12461 15932 12495
rect 15898 12393 15932 12427
rect 15898 12325 15932 12359
rect 15898 12257 15932 12291
rect 15898 12189 15932 12223
rect 15898 12121 15932 12155
rect 15898 12053 15932 12087
rect 15898 11985 15932 12019
rect 15898 11917 15932 11951
rect 15898 11849 15932 11883
rect 15898 11781 15932 11815
rect 15898 11713 15932 11747
rect 15898 11645 15932 11679
rect 15898 11577 15932 11611
rect 15898 11509 15932 11543
rect 15898 11441 15932 11475
rect 15898 11373 15932 11407
rect 15898 11305 15932 11339
rect 15898 11237 15932 11271
rect 15898 11169 15932 11203
rect 15898 11101 15932 11135
rect 15986 13005 16020 13039
rect 15986 12937 16020 12971
rect 15986 12869 16020 12903
rect 15986 12801 16020 12835
rect 15986 12733 16020 12767
rect 15986 12665 16020 12699
rect 15986 12597 16020 12631
rect 15986 12529 16020 12563
rect 15986 12461 16020 12495
rect 15986 12393 16020 12427
rect 15986 12325 16020 12359
rect 15986 12257 16020 12291
rect 15986 12189 16020 12223
rect 15986 12121 16020 12155
rect 15986 12053 16020 12087
rect 15986 11985 16020 12019
rect 15986 11917 16020 11951
rect 15986 11849 16020 11883
rect 15986 11781 16020 11815
rect 15986 11713 16020 11747
rect 15986 11645 16020 11679
rect 15986 11577 16020 11611
rect 15986 11509 16020 11543
rect 15986 11441 16020 11475
rect 15986 11373 16020 11407
rect 15986 11305 16020 11339
rect 15986 11237 16020 11271
rect 15986 11169 16020 11203
rect 15986 11101 16020 11135
rect 16074 13005 16108 13039
rect 16074 12937 16108 12971
rect 16074 12869 16108 12903
rect 16074 12801 16108 12835
rect 16074 12733 16108 12767
rect 16074 12665 16108 12699
rect 16074 12597 16108 12631
rect 16074 12529 16108 12563
rect 16074 12461 16108 12495
rect 16074 12393 16108 12427
rect 16074 12325 16108 12359
rect 16074 12257 16108 12291
rect 16074 12189 16108 12223
rect 16074 12121 16108 12155
rect 16074 12053 16108 12087
rect 16074 11985 16108 12019
rect 16074 11917 16108 11951
rect 16074 11849 16108 11883
rect 16074 11781 16108 11815
rect 16074 11713 16108 11747
rect 16074 11645 16108 11679
rect 16074 11577 16108 11611
rect 16074 11509 16108 11543
rect 16074 11441 16108 11475
rect 16074 11373 16108 11407
rect 16074 11305 16108 11339
rect 16074 11237 16108 11271
rect 16074 11169 16108 11203
rect 16074 11101 16108 11135
rect 16162 13005 16196 13039
rect 16162 12937 16196 12971
rect 16162 12869 16196 12903
rect 16162 12801 16196 12835
rect 16162 12733 16196 12767
rect 16162 12665 16196 12699
rect 16162 12597 16196 12631
rect 16162 12529 16196 12563
rect 16162 12461 16196 12495
rect 16162 12393 16196 12427
rect 16162 12325 16196 12359
rect 16162 12257 16196 12291
rect 16162 12189 16196 12223
rect 16162 12121 16196 12155
rect 16162 12053 16196 12087
rect 16162 11985 16196 12019
rect 16162 11917 16196 11951
rect 16162 11849 16196 11883
rect 16162 11781 16196 11815
rect 16162 11713 16196 11747
rect 16162 11645 16196 11679
rect 16162 11577 16196 11611
rect 16162 11509 16196 11543
rect 16162 11441 16196 11475
rect 16162 11373 16196 11407
rect 16162 11305 16196 11339
rect 16162 11237 16196 11271
rect 16162 11169 16196 11203
rect 16162 11101 16196 11135
rect 16250 13005 16284 13039
rect 16250 12937 16284 12971
rect 16250 12869 16284 12903
rect 16250 12801 16284 12835
rect 16250 12733 16284 12767
rect 16250 12665 16284 12699
rect 16250 12597 16284 12631
rect 16250 12529 16284 12563
rect 16250 12461 16284 12495
rect 16250 12393 16284 12427
rect 16250 12325 16284 12359
rect 16250 12257 16284 12291
rect 16250 12189 16284 12223
rect 16250 12121 16284 12155
rect 16250 12053 16284 12087
rect 16250 11985 16284 12019
rect 16250 11917 16284 11951
rect 16250 11849 16284 11883
rect 16250 11781 16284 11815
rect 16250 11713 16284 11747
rect 16250 11645 16284 11679
rect 16250 11577 16284 11611
rect 16250 11509 16284 11543
rect 16250 11441 16284 11475
rect 16250 11373 16284 11407
rect 16250 11305 16284 11339
rect 16250 11237 16284 11271
rect 16250 11169 16284 11203
rect 16250 11101 16284 11135
rect 16338 13005 16372 13039
rect 16338 12937 16372 12971
rect 16338 12869 16372 12903
rect 16338 12801 16372 12835
rect 16338 12733 16372 12767
rect 16338 12665 16372 12699
rect 16338 12597 16372 12631
rect 16338 12529 16372 12563
rect 16338 12461 16372 12495
rect 16338 12393 16372 12427
rect 16338 12325 16372 12359
rect 16338 12257 16372 12291
rect 16338 12189 16372 12223
rect 16338 12121 16372 12155
rect 16338 12053 16372 12087
rect 16338 11985 16372 12019
rect 16338 11917 16372 11951
rect 16338 11849 16372 11883
rect 16338 11781 16372 11815
rect 16338 11713 16372 11747
rect 16338 11645 16372 11679
rect 16338 11577 16372 11611
rect 16338 11509 16372 11543
rect 16338 11441 16372 11475
rect 16338 11373 16372 11407
rect 16338 11305 16372 11339
rect 16338 11237 16372 11271
rect 16338 11169 16372 11203
rect 16338 11101 16372 11135
rect 16426 13005 16460 13039
rect 16426 12937 16460 12971
rect 16426 12869 16460 12903
rect 16426 12801 16460 12835
rect 16426 12733 16460 12767
rect 16426 12665 16460 12699
rect 16426 12597 16460 12631
rect 16426 12529 16460 12563
rect 16426 12461 16460 12495
rect 16426 12393 16460 12427
rect 16426 12325 16460 12359
rect 16426 12257 16460 12291
rect 16426 12189 16460 12223
rect 16426 12121 16460 12155
rect 16426 12053 16460 12087
rect 16426 11985 16460 12019
rect 16426 11917 16460 11951
rect 16426 11849 16460 11883
rect 16426 11781 16460 11815
rect 16426 11713 16460 11747
rect 16426 11645 16460 11679
rect 16426 11577 16460 11611
rect 16426 11509 16460 11543
rect 16426 11441 16460 11475
rect 16426 11373 16460 11407
rect 16426 11305 16460 11339
rect 16426 11237 16460 11271
rect 16426 11169 16460 11203
rect 16426 11101 16460 11135
rect 16514 13005 16548 13039
rect 16514 12937 16548 12971
rect 16514 12869 16548 12903
rect 16514 12801 16548 12835
rect 16514 12733 16548 12767
rect 16514 12665 16548 12699
rect 16514 12597 16548 12631
rect 16514 12529 16548 12563
rect 16514 12461 16548 12495
rect 16514 12393 16548 12427
rect 16514 12325 16548 12359
rect 16514 12257 16548 12291
rect 16514 12189 16548 12223
rect 16514 12121 16548 12155
rect 16514 12053 16548 12087
rect 16514 11985 16548 12019
rect 16514 11917 16548 11951
rect 16514 11849 16548 11883
rect 16514 11781 16548 11815
rect 16514 11713 16548 11747
rect 16514 11645 16548 11679
rect 16514 11577 16548 11611
rect 16514 11509 16548 11543
rect 16514 11441 16548 11475
rect 16514 11373 16548 11407
rect 16514 11305 16548 11339
rect 16514 11237 16548 11271
rect 16514 11169 16548 11203
rect 16514 11101 16548 11135
rect 16602 13005 16636 13039
rect 16602 12937 16636 12971
rect 16602 12869 16636 12903
rect 16602 12801 16636 12835
rect 16602 12733 16636 12767
rect 16602 12665 16636 12699
rect 16602 12597 16636 12631
rect 16602 12529 16636 12563
rect 16602 12461 16636 12495
rect 16602 12393 16636 12427
rect 16602 12325 16636 12359
rect 16602 12257 16636 12291
rect 16602 12189 16636 12223
rect 16602 12121 16636 12155
rect 16602 12053 16636 12087
rect 16602 11985 16636 12019
rect 16602 11917 16636 11951
rect 16602 11849 16636 11883
rect 16602 11781 16636 11815
rect 16602 11713 16636 11747
rect 16602 11645 16636 11679
rect 16602 11577 16636 11611
rect 16602 11509 16636 11543
rect 16602 11441 16636 11475
rect 16602 11373 16636 11407
rect 16602 11305 16636 11339
rect 16602 11237 16636 11271
rect 16602 11169 16636 11203
rect 16602 11101 16636 11135
rect 16690 13005 16724 13039
rect 16690 12937 16724 12971
rect 16690 12869 16724 12903
rect 16690 12801 16724 12835
rect 16690 12733 16724 12767
rect 16690 12665 16724 12699
rect 16690 12597 16724 12631
rect 16690 12529 16724 12563
rect 16690 12461 16724 12495
rect 16690 12393 16724 12427
rect 16690 12325 16724 12359
rect 16690 12257 16724 12291
rect 16690 12189 16724 12223
rect 16690 12121 16724 12155
rect 16690 12053 16724 12087
rect 16690 11985 16724 12019
rect 16690 11917 16724 11951
rect 16690 11849 16724 11883
rect 16690 11781 16724 11815
rect 16690 11713 16724 11747
rect 16690 11645 16724 11679
rect 16690 11577 16724 11611
rect 16690 11509 16724 11543
rect 16690 11441 16724 11475
rect 16690 11373 16724 11407
rect 16690 11305 16724 11339
rect 16690 11237 16724 11271
rect 16690 11169 16724 11203
rect 16690 11101 16724 11135
rect 16778 13005 16812 13039
rect 16778 12937 16812 12971
rect 16778 12869 16812 12903
rect 16778 12801 16812 12835
rect 16778 12733 16812 12767
rect 16778 12665 16812 12699
rect 16778 12597 16812 12631
rect 16778 12529 16812 12563
rect 16778 12461 16812 12495
rect 16778 12393 16812 12427
rect 16778 12325 16812 12359
rect 16778 12257 16812 12291
rect 16778 12189 16812 12223
rect 16778 12121 16812 12155
rect 16778 12053 16812 12087
rect 16778 11985 16812 12019
rect 16778 11917 16812 11951
rect 16778 11849 16812 11883
rect 16778 11781 16812 11815
rect 16778 11713 16812 11747
rect 16778 11645 16812 11679
rect 16778 11577 16812 11611
rect 16778 11509 16812 11543
rect 16778 11441 16812 11475
rect 16778 11373 16812 11407
rect 16778 11305 16812 11339
rect 16778 11237 16812 11271
rect 16778 11169 16812 11203
rect 16778 11101 16812 11135
rect 16866 13005 16900 13039
rect 16866 12937 16900 12971
rect 16866 12869 16900 12903
rect 16866 12801 16900 12835
rect 16866 12733 16900 12767
rect 16866 12665 16900 12699
rect 16866 12597 16900 12631
rect 16866 12529 16900 12563
rect 16866 12461 16900 12495
rect 16866 12393 16900 12427
rect 16866 12325 16900 12359
rect 16866 12257 16900 12291
rect 16866 12189 16900 12223
rect 16866 12121 16900 12155
rect 16866 12053 16900 12087
rect 16866 11985 16900 12019
rect 16866 11917 16900 11951
rect 16866 11849 16900 11883
rect 16866 11781 16900 11815
rect 16866 11713 16900 11747
rect 16866 11645 16900 11679
rect 16866 11577 16900 11611
rect 16866 11509 16900 11543
rect 16866 11441 16900 11475
rect 16866 11373 16900 11407
rect 16866 11305 16900 11339
rect 16866 11237 16900 11271
rect 16866 11169 16900 11203
rect 16866 11101 16900 11135
rect 16954 13005 16988 13039
rect 16954 12937 16988 12971
rect 16954 12869 16988 12903
rect 16954 12801 16988 12835
rect 16954 12733 16988 12767
rect 16954 12665 16988 12699
rect 16954 12597 16988 12631
rect 16954 12529 16988 12563
rect 16954 12461 16988 12495
rect 16954 12393 16988 12427
rect 16954 12325 16988 12359
rect 16954 12257 16988 12291
rect 16954 12189 16988 12223
rect 16954 12121 16988 12155
rect 16954 12053 16988 12087
rect 16954 11985 16988 12019
rect 16954 11917 16988 11951
rect 16954 11849 16988 11883
rect 16954 11781 16988 11815
rect 16954 11713 16988 11747
rect 16954 11645 16988 11679
rect 16954 11577 16988 11611
rect 16954 11509 16988 11543
rect 16954 11441 16988 11475
rect 16954 11373 16988 11407
rect 16954 11305 16988 11339
rect 16954 11237 16988 11271
rect 16954 11169 16988 11203
rect 16954 11101 16988 11135
rect 17042 13005 17076 13039
rect 17042 12937 17076 12971
rect 17042 12869 17076 12903
rect 17042 12801 17076 12835
rect 17042 12733 17076 12767
rect 17042 12665 17076 12699
rect 17042 12597 17076 12631
rect 17042 12529 17076 12563
rect 17042 12461 17076 12495
rect 17042 12393 17076 12427
rect 17042 12325 17076 12359
rect 17042 12257 17076 12291
rect 17042 12189 17076 12223
rect 17042 12121 17076 12155
rect 17042 12053 17076 12087
rect 17042 11985 17076 12019
rect 17042 11917 17076 11951
rect 17042 11849 17076 11883
rect 17042 11781 17076 11815
rect 17042 11713 17076 11747
rect 17042 11645 17076 11679
rect 17042 11577 17076 11611
rect 17042 11509 17076 11543
rect 17042 11441 17076 11475
rect 17042 11373 17076 11407
rect 17042 11305 17076 11339
rect 17042 11237 17076 11271
rect 17042 11169 17076 11203
rect 17042 11101 17076 11135
rect 17130 13005 17164 13039
rect 17130 12937 17164 12971
rect 17130 12869 17164 12903
rect 17130 12801 17164 12835
rect 17130 12733 17164 12767
rect 17130 12665 17164 12699
rect 17130 12597 17164 12631
rect 17130 12529 17164 12563
rect 17130 12461 17164 12495
rect 17130 12393 17164 12427
rect 17130 12325 17164 12359
rect 17130 12257 17164 12291
rect 17130 12189 17164 12223
rect 17130 12121 17164 12155
rect 17130 12053 17164 12087
rect 17130 11985 17164 12019
rect 17130 11917 17164 11951
rect 17130 11849 17164 11883
rect 17130 11781 17164 11815
rect 17130 11713 17164 11747
rect 17130 11645 17164 11679
rect 17130 11577 17164 11611
rect 17130 11509 17164 11543
rect 17130 11441 17164 11475
rect 17130 11373 17164 11407
rect 17130 11305 17164 11339
rect 17130 11237 17164 11271
rect 17130 11169 17164 11203
rect 17130 11101 17164 11135
rect 17218 13005 17252 13039
rect 17218 12937 17252 12971
rect 17218 12869 17252 12903
rect 17218 12801 17252 12835
rect 17218 12733 17252 12767
rect 17218 12665 17252 12699
rect 17218 12597 17252 12631
rect 17218 12529 17252 12563
rect 17218 12461 17252 12495
rect 17218 12393 17252 12427
rect 17218 12325 17252 12359
rect 17218 12257 17252 12291
rect 17218 12189 17252 12223
rect 17218 12121 17252 12155
rect 17218 12053 17252 12087
rect 17218 11985 17252 12019
rect 17218 11917 17252 11951
rect 17218 11849 17252 11883
rect 17218 11781 17252 11815
rect 17218 11713 17252 11747
rect 17218 11645 17252 11679
rect 17218 11577 17252 11611
rect 17218 11509 17252 11543
rect 17218 11441 17252 11475
rect 17218 11373 17252 11407
rect 17218 11305 17252 11339
rect 17218 11237 17252 11271
rect 17218 11169 17252 11203
rect 17218 11101 17252 11135
rect 17306 13005 17340 13039
rect 17306 12937 17340 12971
rect 17306 12869 17340 12903
rect 17306 12801 17340 12835
rect 17306 12733 17340 12767
rect 17306 12665 17340 12699
rect 17306 12597 17340 12631
rect 17306 12529 17340 12563
rect 17306 12461 17340 12495
rect 17306 12393 17340 12427
rect 17306 12325 17340 12359
rect 17306 12257 17340 12291
rect 17306 12189 17340 12223
rect 17306 12121 17340 12155
rect 17306 12053 17340 12087
rect 17306 11985 17340 12019
rect 17306 11917 17340 11951
rect 17306 11849 17340 11883
rect 17306 11781 17340 11815
rect 17306 11713 17340 11747
rect 17306 11645 17340 11679
rect 17306 11577 17340 11611
rect 17306 11509 17340 11543
rect 17306 11441 17340 11475
rect 17306 11373 17340 11407
rect 17306 11305 17340 11339
rect 17306 11237 17340 11271
rect 17306 11169 17340 11203
rect 17306 11101 17340 11135
rect 17394 13005 17428 13039
rect 17394 12937 17428 12971
rect 17394 12869 17428 12903
rect 17394 12801 17428 12835
rect 17394 12733 17428 12767
rect 17394 12665 17428 12699
rect 17394 12597 17428 12631
rect 17394 12529 17428 12563
rect 17394 12461 17428 12495
rect 17394 12393 17428 12427
rect 17394 12325 17428 12359
rect 17394 12257 17428 12291
rect 17394 12189 17428 12223
rect 17394 12121 17428 12155
rect 17394 12053 17428 12087
rect 17394 11985 17428 12019
rect 17394 11917 17428 11951
rect 17394 11849 17428 11883
rect 17394 11781 17428 11815
rect 17394 11713 17428 11747
rect 17394 11645 17428 11679
rect 17394 11577 17428 11611
rect 17394 11509 17428 11543
rect 17394 11441 17428 11475
rect 17394 11373 17428 11407
rect 17394 11305 17428 11339
rect 17394 11237 17428 11271
rect 17394 11169 17428 11203
rect 17394 11101 17428 11135
rect 17482 13005 17516 13039
rect 17482 12937 17516 12971
rect 17482 12869 17516 12903
rect 17482 12801 17516 12835
rect 17482 12733 17516 12767
rect 17482 12665 17516 12699
rect 17482 12597 17516 12631
rect 17482 12529 17516 12563
rect 17482 12461 17516 12495
rect 17482 12393 17516 12427
rect 17482 12325 17516 12359
rect 17482 12257 17516 12291
rect 17482 12189 17516 12223
rect 17482 12121 17516 12155
rect 17482 12053 17516 12087
rect 17482 11985 17516 12019
rect 17482 11917 17516 11951
rect 17482 11849 17516 11883
rect 17482 11781 17516 11815
rect 17482 11713 17516 11747
rect 17482 11645 17516 11679
rect 17482 11577 17516 11611
rect 17482 11509 17516 11543
rect 17482 11441 17516 11475
rect 17482 11373 17516 11407
rect 17482 11305 17516 11339
rect 17482 11237 17516 11271
rect 17482 11169 17516 11203
rect 17482 11101 17516 11135
<< pdiffc >>
rect 15830 23124 15864 23158
rect 15830 23056 15864 23090
rect 15830 22988 15864 23022
rect 15830 22920 15864 22954
rect 15830 22852 15864 22886
rect 15830 22784 15864 22818
rect 15830 22716 15864 22750
rect 15830 22648 15864 22682
rect 15830 22580 15864 22614
rect 15830 22512 15864 22546
rect 15830 22444 15864 22478
rect 15830 22376 15864 22410
rect 15830 22308 15864 22342
rect 15830 22240 15864 22274
rect 15830 22172 15864 22206
rect 15830 22104 15864 22138
rect 15830 22036 15864 22070
rect 15830 21968 15864 22002
rect 15830 21900 15864 21934
rect 15830 21832 15864 21866
rect 15830 21764 15864 21798
rect 15830 21696 15864 21730
rect 15830 21628 15864 21662
rect 15830 21560 15864 21594
rect 15830 21492 15864 21526
rect 15830 21424 15864 21458
rect 15830 21356 15864 21390
rect 15830 21288 15864 21322
rect 15830 21220 15864 21254
rect 15926 23124 15960 23158
rect 15926 23056 15960 23090
rect 15926 22988 15960 23022
rect 15926 22920 15960 22954
rect 15926 22852 15960 22886
rect 15926 22784 15960 22818
rect 15926 22716 15960 22750
rect 15926 22648 15960 22682
rect 15926 22580 15960 22614
rect 15926 22512 15960 22546
rect 15926 22444 15960 22478
rect 15926 22376 15960 22410
rect 15926 22308 15960 22342
rect 15926 22240 15960 22274
rect 15926 22172 15960 22206
rect 15926 22104 15960 22138
rect 15926 22036 15960 22070
rect 15926 21968 15960 22002
rect 15926 21900 15960 21934
rect 15926 21832 15960 21866
rect 15926 21764 15960 21798
rect 15926 21696 15960 21730
rect 15926 21628 15960 21662
rect 15926 21560 15960 21594
rect 15926 21492 15960 21526
rect 15926 21424 15960 21458
rect 15926 21356 15960 21390
rect 15926 21288 15960 21322
rect 15926 21220 15960 21254
rect 16022 23124 16056 23158
rect 16022 23056 16056 23090
rect 16022 22988 16056 23022
rect 16022 22920 16056 22954
rect 16022 22852 16056 22886
rect 16022 22784 16056 22818
rect 16022 22716 16056 22750
rect 16022 22648 16056 22682
rect 16022 22580 16056 22614
rect 16022 22512 16056 22546
rect 16022 22444 16056 22478
rect 16022 22376 16056 22410
rect 16022 22308 16056 22342
rect 16022 22240 16056 22274
rect 16022 22172 16056 22206
rect 16022 22104 16056 22138
rect 16022 22036 16056 22070
rect 16022 21968 16056 22002
rect 16022 21900 16056 21934
rect 16022 21832 16056 21866
rect 16022 21764 16056 21798
rect 16022 21696 16056 21730
rect 16022 21628 16056 21662
rect 16022 21560 16056 21594
rect 16022 21492 16056 21526
rect 16022 21424 16056 21458
rect 16022 21356 16056 21390
rect 16022 21288 16056 21322
rect 16022 21220 16056 21254
rect 16118 23124 16152 23158
rect 16118 23056 16152 23090
rect 16118 22988 16152 23022
rect 16118 22920 16152 22954
rect 16118 22852 16152 22886
rect 16118 22784 16152 22818
rect 16118 22716 16152 22750
rect 16118 22648 16152 22682
rect 16118 22580 16152 22614
rect 16118 22512 16152 22546
rect 16118 22444 16152 22478
rect 16118 22376 16152 22410
rect 16118 22308 16152 22342
rect 16118 22240 16152 22274
rect 16118 22172 16152 22206
rect 16118 22104 16152 22138
rect 16118 22036 16152 22070
rect 16118 21968 16152 22002
rect 16118 21900 16152 21934
rect 16118 21832 16152 21866
rect 16118 21764 16152 21798
rect 16118 21696 16152 21730
rect 16118 21628 16152 21662
rect 16118 21560 16152 21594
rect 16118 21492 16152 21526
rect 16118 21424 16152 21458
rect 16118 21356 16152 21390
rect 16118 21288 16152 21322
rect 16118 21220 16152 21254
rect 17092 15878 17126 15912
rect 17092 15810 17126 15844
rect 17092 15742 17126 15776
rect 17092 15674 17126 15708
rect 17092 15606 17126 15640
rect 17092 15538 17126 15572
rect 17092 15470 17126 15504
rect 17092 15402 17126 15436
rect 17092 15334 17126 15368
rect 17092 15266 17126 15300
rect 17092 15198 17126 15232
rect 17092 15130 17126 15164
rect 17092 15062 17126 15096
rect 17092 14994 17126 15028
rect 17092 14926 17126 14960
rect 17092 14858 17126 14892
rect 17092 14790 17126 14824
rect 17092 14722 17126 14756
rect 17092 14654 17126 14688
rect 17092 14586 17126 14620
rect 17092 14518 17126 14552
rect 17092 14450 17126 14484
rect 17092 14382 17126 14416
rect 17092 14314 17126 14348
rect 17092 14246 17126 14280
rect 17092 14178 17126 14212
rect 17092 14110 17126 14144
rect 17092 14042 17126 14076
rect 17092 13974 17126 14008
rect 17188 15878 17222 15912
rect 17188 15810 17222 15844
rect 17188 15742 17222 15776
rect 17188 15674 17222 15708
rect 17188 15606 17222 15640
rect 17188 15538 17222 15572
rect 17188 15470 17222 15504
rect 17188 15402 17222 15436
rect 17188 15334 17222 15368
rect 17188 15266 17222 15300
rect 17188 15198 17222 15232
rect 17188 15130 17222 15164
rect 17188 15062 17222 15096
rect 17188 14994 17222 15028
rect 17188 14926 17222 14960
rect 17188 14858 17222 14892
rect 17188 14790 17222 14824
rect 17188 14722 17222 14756
rect 17188 14654 17222 14688
rect 17188 14586 17222 14620
rect 17188 14518 17222 14552
rect 17188 14450 17222 14484
rect 17188 14382 17222 14416
rect 17188 14314 17222 14348
rect 17188 14246 17222 14280
rect 17188 14178 17222 14212
rect 17188 14110 17222 14144
rect 17188 14042 17222 14076
rect 17188 13974 17222 14008
rect 17284 15878 17318 15912
rect 17284 15810 17318 15844
rect 17284 15742 17318 15776
rect 17284 15674 17318 15708
rect 17284 15606 17318 15640
rect 17284 15538 17318 15572
rect 17284 15470 17318 15504
rect 17284 15402 17318 15436
rect 17284 15334 17318 15368
rect 17284 15266 17318 15300
rect 17284 15198 17318 15232
rect 17284 15130 17318 15164
rect 17284 15062 17318 15096
rect 17284 14994 17318 15028
rect 17284 14926 17318 14960
rect 17284 14858 17318 14892
rect 17284 14790 17318 14824
rect 17284 14722 17318 14756
rect 17284 14654 17318 14688
rect 17284 14586 17318 14620
rect 17284 14518 17318 14552
rect 17284 14450 17318 14484
rect 17284 14382 17318 14416
rect 17284 14314 17318 14348
rect 17284 14246 17318 14280
rect 17284 14178 17318 14212
rect 17284 14110 17318 14144
rect 17284 14042 17318 14076
rect 17284 13974 17318 14008
rect 17380 15878 17414 15912
rect 17380 15810 17414 15844
rect 17380 15742 17414 15776
rect 17380 15674 17414 15708
rect 17380 15606 17414 15640
rect 17380 15538 17414 15572
rect 17380 15470 17414 15504
rect 17380 15402 17414 15436
rect 17380 15334 17414 15368
rect 17380 15266 17414 15300
rect 17380 15198 17414 15232
rect 17380 15130 17414 15164
rect 17380 15062 17414 15096
rect 17380 14994 17414 15028
rect 17380 14926 17414 14960
rect 17380 14858 17414 14892
rect 17380 14790 17414 14824
rect 17380 14722 17414 14756
rect 17380 14654 17414 14688
rect 17380 14586 17414 14620
rect 17380 14518 17414 14552
rect 17380 14450 17414 14484
rect 17380 14382 17414 14416
rect 17380 14314 17414 14348
rect 17380 14246 17414 14280
rect 17380 14178 17414 14212
rect 17380 14110 17414 14144
rect 17380 14042 17414 14076
rect 17380 13974 17414 14008
<< psubdiff >>
rect 12916 24712 13023 24746
rect 13057 24712 13091 24746
rect 13125 24712 13159 24746
rect 13193 24712 13227 24746
rect 13261 24712 13295 24746
rect 13329 24712 13363 24746
rect 13397 24712 13431 24746
rect 13465 24712 13499 24746
rect 13533 24712 13567 24746
rect 13601 24712 13635 24746
rect 13669 24712 13703 24746
rect 13737 24712 13771 24746
rect 13805 24712 13839 24746
rect 13873 24712 13907 24746
rect 13941 24712 13975 24746
rect 14009 24712 14043 24746
rect 14077 24712 14111 24746
rect 14145 24712 14179 24746
rect 14213 24712 14247 24746
rect 14281 24712 14315 24746
rect 14349 24712 14383 24746
rect 14417 24712 14451 24746
rect 14485 24712 14519 24746
rect 14553 24712 14587 24746
rect 14621 24712 14655 24746
rect 14689 24712 14723 24746
rect 14757 24712 14791 24746
rect 14825 24712 14859 24746
rect 14893 24712 14927 24746
rect 14961 24712 14995 24746
rect 15029 24712 15063 24746
rect 15097 24712 15131 24746
rect 15165 24712 15199 24746
rect 15233 24712 15267 24746
rect 15301 24712 15335 24746
rect 15369 24712 15403 24746
rect 15437 24712 15471 24746
rect 15505 24712 15539 24746
rect 15573 24712 15607 24746
rect 15641 24712 15675 24746
rect 15709 24712 15743 24746
rect 15777 24712 15811 24746
rect 15845 24712 15879 24746
rect 15913 24712 15947 24746
rect 15981 24712 16015 24746
rect 16049 24712 16083 24746
rect 16117 24712 16151 24746
rect 16185 24712 16219 24746
rect 16253 24712 16287 24746
rect 16321 24712 16355 24746
rect 16389 24712 16423 24746
rect 16457 24712 16491 24746
rect 16525 24712 16559 24746
rect 16593 24712 16627 24746
rect 16661 24712 16695 24746
rect 16729 24712 16763 24746
rect 16797 24712 16831 24746
rect 16865 24712 16899 24746
rect 16933 24712 17040 24746
rect 12916 24632 12950 24712
rect 17006 24632 17040 24712
rect 12916 24564 12950 24598
rect 17006 24564 17040 24598
rect 12916 24450 12950 24530
rect 17006 24450 17040 24530
rect 12916 24416 13023 24450
rect 13057 24416 13091 24450
rect 13125 24416 13159 24450
rect 13193 24416 13227 24450
rect 13261 24416 13295 24450
rect 13329 24416 13363 24450
rect 13397 24416 13431 24450
rect 13465 24416 13499 24450
rect 13533 24416 13567 24450
rect 13601 24416 13635 24450
rect 13669 24416 13703 24450
rect 13737 24416 13771 24450
rect 13805 24416 13839 24450
rect 13873 24416 13907 24450
rect 13941 24416 13975 24450
rect 14009 24416 14043 24450
rect 14077 24416 14111 24450
rect 14145 24416 14179 24450
rect 14213 24416 14247 24450
rect 14281 24416 14315 24450
rect 14349 24416 14383 24450
rect 14417 24416 14451 24450
rect 14485 24416 14519 24450
rect 14553 24416 14587 24450
rect 14621 24416 14655 24450
rect 14689 24416 14723 24450
rect 14757 24416 14791 24450
rect 14825 24416 14859 24450
rect 14893 24416 14927 24450
rect 14961 24416 14995 24450
rect 15029 24416 15063 24450
rect 15097 24416 15131 24450
rect 15165 24416 15199 24450
rect 15233 24416 15267 24450
rect 15301 24416 15335 24450
rect 15369 24416 15403 24450
rect 15437 24416 15471 24450
rect 15505 24416 15539 24450
rect 15573 24416 15607 24450
rect 15641 24416 15675 24450
rect 15709 24416 15743 24450
rect 15777 24416 15811 24450
rect 15845 24416 15879 24450
rect 15913 24416 15947 24450
rect 15981 24416 16015 24450
rect 16049 24416 16083 24450
rect 16117 24416 16151 24450
rect 16185 24416 16219 24450
rect 16253 24416 16287 24450
rect 16321 24416 16355 24450
rect 16389 24416 16423 24450
rect 16457 24416 16491 24450
rect 16525 24416 16559 24450
rect 16593 24416 16627 24450
rect 16661 24416 16695 24450
rect 16729 24416 16763 24450
rect 16797 24416 16831 24450
rect 16865 24416 16899 24450
rect 16933 24416 17040 24450
rect 16548 24180 16666 24214
rect 16700 24180 16734 24214
rect 16768 24180 16802 24214
rect 16836 24180 16870 24214
rect 16904 24180 16938 24214
rect 16972 24180 17006 24214
rect 17040 24180 17074 24214
rect 17108 24180 17142 24214
rect 17176 24180 17210 24214
rect 17244 24180 17278 24214
rect 17312 24180 17346 24214
rect 17380 24180 17414 24214
rect 17448 24180 17482 24214
rect 17516 24180 17550 24214
rect 17584 24180 17618 24214
rect 17652 24180 17770 24214
rect 16548 24111 16582 24180
rect 12946 24032 13075 24066
rect 13109 24032 13143 24066
rect 13177 24032 13211 24066
rect 13245 24032 13279 24066
rect 13313 24032 13347 24066
rect 13381 24032 13415 24066
rect 13449 24032 13483 24066
rect 13517 24032 13551 24066
rect 13585 24032 13619 24066
rect 13653 24032 13687 24066
rect 13721 24032 13755 24066
rect 13789 24032 13823 24066
rect 13857 24032 13891 24066
rect 13925 24032 13959 24066
rect 13993 24032 14027 24066
rect 14061 24032 14095 24066
rect 14129 24032 14163 24066
rect 14197 24032 14231 24066
rect 14265 24032 14299 24066
rect 14333 24032 14367 24066
rect 14401 24032 14435 24066
rect 14469 24032 14503 24066
rect 14537 24032 14571 24066
rect 14605 24032 14639 24066
rect 14673 24032 14707 24066
rect 14741 24032 14870 24066
rect 12946 23952 12980 24032
rect 14836 23952 14870 24032
rect 12946 23884 12980 23918
rect 14836 23884 14870 23918
rect 12946 23770 12980 23850
rect 14836 23770 14870 23850
rect 12946 23736 13075 23770
rect 13109 23736 13143 23770
rect 13177 23736 13211 23770
rect 13245 23736 13279 23770
rect 13313 23736 13347 23770
rect 13381 23736 13415 23770
rect 13449 23736 13483 23770
rect 13517 23736 13551 23770
rect 13585 23736 13619 23770
rect 13653 23736 13687 23770
rect 13721 23736 13755 23770
rect 13789 23736 13823 23770
rect 13857 23736 13891 23770
rect 13925 23736 13959 23770
rect 13993 23736 14027 23770
rect 14061 23736 14095 23770
rect 14129 23736 14163 23770
rect 14197 23736 14231 23770
rect 14265 23736 14299 23770
rect 14333 23736 14367 23770
rect 14401 23736 14435 23770
rect 14469 23736 14503 23770
rect 14537 23736 14571 23770
rect 14605 23736 14639 23770
rect 14673 23736 14707 23770
rect 14741 23736 14870 23770
rect 16548 24043 16582 24077
rect 17736 24111 17770 24180
rect 17736 24043 17770 24077
rect 16548 23975 16582 24009
rect 16548 23907 16582 23941
rect 16548 23839 16582 23873
rect 16548 23771 16582 23805
rect 16548 23703 16582 23737
rect 16548 23635 16582 23669
rect 16548 23567 16582 23601
rect 16548 23499 16582 23533
rect 16548 23431 16582 23465
rect 15176 23326 15290 23360
rect 15324 23326 15358 23360
rect 15392 23326 15506 23360
rect 13856 23290 13980 23324
rect 14014 23290 14048 23324
rect 14082 23290 14116 23324
rect 14150 23290 14184 23324
rect 14218 23290 14252 23324
rect 14286 23290 14320 23324
rect 14354 23290 14388 23324
rect 14422 23290 14456 23324
rect 14490 23290 14524 23324
rect 14558 23290 14592 23324
rect 14626 23290 14660 23324
rect 14694 23290 14728 23324
rect 14762 23290 14886 23324
rect 13856 23221 13890 23290
rect 13856 23153 13890 23187
rect 14852 23221 14886 23290
rect 14852 23153 14886 23187
rect 13856 23085 13890 23119
rect 13856 23017 13890 23051
rect 13856 22949 13890 22983
rect 13856 22881 13890 22915
rect 13856 22813 13890 22847
rect 13856 22745 13890 22779
rect 13856 22677 13890 22711
rect 13856 22609 13890 22643
rect 13856 22541 13890 22575
rect 13856 22473 13890 22507
rect 13856 22405 13890 22439
rect 13856 22337 13890 22371
rect 13856 22269 13890 22303
rect 13856 22201 13890 22235
rect 13356 22166 13470 22200
rect 13504 22166 13538 22200
rect 13572 22166 13686 22200
rect 13356 22081 13390 22166
rect 13652 22081 13686 22166
rect 13356 22013 13390 22047
rect 13356 21945 13390 21979
rect 13356 21877 13390 21911
rect 13356 21809 13390 21843
rect 13356 21741 13390 21775
rect 13356 21673 13390 21707
rect 13356 21605 13390 21639
rect 13356 21537 13390 21571
rect 13356 21469 13390 21503
rect 13356 21401 13390 21435
rect 13356 21333 13390 21367
rect 13356 21265 13390 21299
rect 13356 21197 13390 21231
rect 13356 21129 13390 21163
rect 13652 22013 13686 22047
rect 13652 21945 13686 21979
rect 13652 21877 13686 21911
rect 13652 21809 13686 21843
rect 13652 21741 13686 21775
rect 13652 21673 13686 21707
rect 13652 21605 13686 21639
rect 13652 21537 13686 21571
rect 13652 21469 13686 21503
rect 13652 21401 13686 21435
rect 13652 21333 13686 21367
rect 13652 21265 13686 21299
rect 13652 21197 13686 21231
rect 13652 21129 13686 21163
rect 13356 21010 13390 21095
rect 13652 21010 13686 21095
rect 13356 20976 13470 21010
rect 13504 20976 13538 21010
rect 13572 20976 13686 21010
rect 13856 22133 13890 22167
rect 13856 22065 13890 22099
rect 13856 21997 13890 22031
rect 13856 21929 13890 21963
rect 13856 21861 13890 21895
rect 13856 21793 13890 21827
rect 13856 21725 13890 21759
rect 13856 21657 13890 21691
rect 13856 21589 13890 21623
rect 13856 21521 13890 21555
rect 13856 21453 13890 21487
rect 13856 21385 13890 21419
rect 13856 21317 13890 21351
rect 13856 21249 13890 21283
rect 13856 21181 13890 21215
rect 14852 23085 14886 23119
rect 14852 23017 14886 23051
rect 14852 22949 14886 22983
rect 14852 22881 14886 22915
rect 14852 22813 14886 22847
rect 14852 22745 14886 22779
rect 14852 22677 14886 22711
rect 14852 22609 14886 22643
rect 14852 22541 14886 22575
rect 14852 22473 14886 22507
rect 14852 22405 14886 22439
rect 14852 22337 14886 22371
rect 14852 22269 14886 22303
rect 14852 22201 14886 22235
rect 14852 22133 14886 22167
rect 14852 22065 14886 22099
rect 14852 21997 14886 22031
rect 14852 21929 14886 21963
rect 14852 21861 14886 21895
rect 14852 21793 14886 21827
rect 14852 21725 14886 21759
rect 14852 21657 14886 21691
rect 14852 21589 14886 21623
rect 14852 21521 14886 21555
rect 14852 21453 14886 21487
rect 14852 21385 14886 21419
rect 14852 21317 14886 21351
rect 14852 21249 14886 21283
rect 14852 21181 14886 21215
rect 13856 21113 13890 21147
rect 13856 21010 13890 21079
rect 14852 21113 14886 21147
rect 14852 21010 14886 21079
rect 13856 20976 13980 21010
rect 14014 20976 14048 21010
rect 14082 20976 14116 21010
rect 14150 20976 14184 21010
rect 14218 20976 14252 21010
rect 14286 20976 14320 21010
rect 14354 20976 14388 21010
rect 14422 20976 14456 21010
rect 14490 20976 14524 21010
rect 14558 20976 14592 21010
rect 14626 20976 14660 21010
rect 14694 20976 14728 21010
rect 14762 20976 14886 21010
rect 15176 23249 15210 23326
rect 15472 23249 15506 23326
rect 15176 23181 15210 23215
rect 15176 23113 15210 23147
rect 15176 23045 15210 23079
rect 15176 22977 15210 23011
rect 15176 22909 15210 22943
rect 15176 22841 15210 22875
rect 15176 22773 15210 22807
rect 15176 22705 15210 22739
rect 15176 22637 15210 22671
rect 15176 22569 15210 22603
rect 15176 22501 15210 22535
rect 15176 22433 15210 22467
rect 15176 22365 15210 22399
rect 15176 22297 15210 22331
rect 15176 22229 15210 22263
rect 15176 22161 15210 22195
rect 15176 22093 15210 22127
rect 15176 22025 15210 22059
rect 15176 21957 15210 21991
rect 15176 21889 15210 21923
rect 15176 21821 15210 21855
rect 15176 21753 15210 21787
rect 15176 21685 15210 21719
rect 15176 21617 15210 21651
rect 15176 21549 15210 21583
rect 15176 21481 15210 21515
rect 15176 21413 15210 21447
rect 15176 21345 15210 21379
rect 15176 21277 15210 21311
rect 15176 21209 15210 21243
rect 15176 21141 15210 21175
rect 15472 23181 15506 23215
rect 15472 23113 15506 23147
rect 15472 23045 15506 23079
rect 15472 22977 15506 23011
rect 15472 22909 15506 22943
rect 15472 22841 15506 22875
rect 15472 22773 15506 22807
rect 15472 22705 15506 22739
rect 15472 22637 15506 22671
rect 15472 22569 15506 22603
rect 15472 22501 15506 22535
rect 15472 22433 15506 22467
rect 15472 22365 15506 22399
rect 15472 22297 15506 22331
rect 15472 22229 15506 22263
rect 15472 22161 15506 22195
rect 15472 22093 15506 22127
rect 15472 22025 15506 22059
rect 15472 21957 15506 21991
rect 15472 21889 15506 21923
rect 15472 21821 15506 21855
rect 15472 21753 15506 21787
rect 15472 21685 15506 21719
rect 15472 21617 15506 21651
rect 15472 21549 15506 21583
rect 15472 21481 15506 21515
rect 15472 21413 15506 21447
rect 15472 21345 15506 21379
rect 15472 21277 15506 21311
rect 15472 21209 15506 21243
rect 15472 21141 15506 21175
rect 15176 21030 15210 21107
rect 15472 21030 15506 21107
rect 15176 20996 15290 21030
rect 15324 20996 15358 21030
rect 15392 20996 15506 21030
rect 16548 23363 16582 23397
rect 16548 23295 16582 23329
rect 16548 23227 16582 23261
rect 16548 23159 16582 23193
rect 16548 23091 16582 23125
rect 16548 23023 16582 23057
rect 16548 22955 16582 22989
rect 16548 22887 16582 22921
rect 16548 22819 16582 22853
rect 16548 22751 16582 22785
rect 16548 22683 16582 22717
rect 16548 22615 16582 22649
rect 16548 22547 16582 22581
rect 16548 22479 16582 22513
rect 16548 22411 16582 22445
rect 16548 22343 16582 22377
rect 16548 22275 16582 22309
rect 16548 22207 16582 22241
rect 16548 22139 16582 22173
rect 16548 22071 16582 22105
rect 17736 23975 17770 24009
rect 17736 23907 17770 23941
rect 17736 23839 17770 23873
rect 17736 23771 17770 23805
rect 17736 23703 17770 23737
rect 17736 23635 17770 23669
rect 17736 23567 17770 23601
rect 17736 23499 17770 23533
rect 17736 23431 17770 23465
rect 17736 23363 17770 23397
rect 17736 23295 17770 23329
rect 17736 23227 17770 23261
rect 17736 23159 17770 23193
rect 17736 23091 17770 23125
rect 17736 23023 17770 23057
rect 17736 22955 17770 22989
rect 17736 22887 17770 22921
rect 17736 22819 17770 22853
rect 17736 22751 17770 22785
rect 17736 22683 17770 22717
rect 17736 22615 17770 22649
rect 17736 22547 17770 22581
rect 17736 22479 17770 22513
rect 17736 22411 17770 22445
rect 17736 22343 17770 22377
rect 17736 22275 17770 22309
rect 17736 22207 17770 22241
rect 17736 22139 17770 22173
rect 17736 22071 17770 22105
rect 16548 22003 16582 22037
rect 16548 21900 16582 21969
rect 17736 22003 17770 22037
rect 17736 21900 17770 21969
rect 16548 21866 16666 21900
rect 16700 21866 16734 21900
rect 16768 21866 16802 21900
rect 16836 21866 16870 21900
rect 16904 21866 16938 21900
rect 16972 21866 17006 21900
rect 17040 21866 17074 21900
rect 17108 21866 17142 21900
rect 17176 21866 17210 21900
rect 17244 21866 17278 21900
rect 17312 21866 17346 21900
rect 17380 21866 17414 21900
rect 17448 21866 17482 21900
rect 17516 21866 17550 21900
rect 17584 21866 17618 21900
rect 17652 21866 17770 21900
rect 16656 21446 16770 21480
rect 16804 21446 16838 21480
rect 16872 21446 16986 21480
rect 16656 21359 16690 21446
rect 16952 21359 16986 21446
rect 16656 21291 16690 21325
rect 16656 21223 16690 21257
rect 16656 21155 16690 21189
rect 16656 21087 16690 21121
rect 16656 21019 16690 21053
rect 16656 20951 16690 20985
rect 16656 20883 16690 20917
rect 16656 20815 16690 20849
rect 16656 20747 16690 20781
rect 16656 20679 16690 20713
rect 14716 20586 14826 20620
rect 14860 20586 14894 20620
rect 14928 20586 14962 20620
rect 14996 20586 15030 20620
rect 15064 20586 15098 20620
rect 15132 20586 15166 20620
rect 15200 20586 15234 20620
rect 15268 20586 15302 20620
rect 15336 20586 15370 20620
rect 15404 20586 15438 20620
rect 15472 20586 15506 20620
rect 15540 20586 15650 20620
rect 14716 20500 14750 20586
rect 14716 20432 14750 20466
rect 15616 20500 15650 20586
rect 14716 20364 14750 20398
rect 14716 20296 14750 20330
rect 14716 20228 14750 20262
rect 14716 20160 14750 20194
rect 14716 20092 14750 20126
rect 14716 20024 14750 20058
rect 14716 19956 14750 19990
rect 14716 19888 14750 19922
rect 13182 19826 13286 19860
rect 13320 19826 13354 19860
rect 13388 19826 13422 19860
rect 13456 19826 13490 19860
rect 13524 19826 13558 19860
rect 13592 19826 13626 19860
rect 13660 19826 13694 19860
rect 13728 19826 13762 19860
rect 13796 19826 13830 19860
rect 13864 19826 13898 19860
rect 13932 19826 13966 19860
rect 14000 19826 14034 19860
rect 14068 19826 14102 19860
rect 14136 19826 14170 19860
rect 14204 19826 14238 19860
rect 14272 19826 14306 19860
rect 14340 19826 14444 19860
rect 13182 19755 13216 19826
rect 14410 19755 14444 19826
rect 13182 19687 13216 19721
rect 13182 19619 13216 19653
rect 14410 19687 14444 19721
rect 14410 19619 14444 19653
rect 13182 19551 13216 19585
rect 13182 19483 13216 19517
rect 13182 19415 13216 19449
rect 13182 19347 13216 19381
rect 14410 19551 14444 19585
rect 14410 19483 14444 19517
rect 14410 19415 14444 19449
rect 14410 19347 14444 19381
rect 13182 19279 13216 19313
rect 13182 19211 13216 19245
rect 14410 19279 14444 19313
rect 14410 19211 14444 19245
rect 13182 19143 13216 19177
rect 13182 19075 13216 19109
rect 13182 19007 13216 19041
rect 13182 18939 13216 18973
rect 14410 19143 14444 19177
rect 14410 19075 14444 19109
rect 14410 19007 14444 19041
rect 14716 19820 14750 19854
rect 14716 19752 14750 19786
rect 14716 19684 14750 19718
rect 14716 19616 14750 19650
rect 14716 19548 14750 19582
rect 14716 19480 14750 19514
rect 14716 19412 14750 19446
rect 14716 19344 14750 19378
rect 14716 19276 14750 19310
rect 14716 19208 14750 19242
rect 14716 19140 14750 19174
rect 15616 20432 15650 20466
rect 15616 20364 15650 20398
rect 15616 20296 15650 20330
rect 15616 20228 15650 20262
rect 15616 20160 15650 20194
rect 16656 20611 16690 20645
rect 16656 20543 16690 20577
rect 16656 20475 16690 20509
rect 16656 20407 16690 20441
rect 16656 20339 16690 20373
rect 16656 20271 16690 20305
rect 16656 20203 16690 20237
rect 16656 20135 16690 20169
rect 15616 20092 15650 20126
rect 15616 20024 15650 20058
rect 15616 19956 15650 19990
rect 15616 19888 15650 19922
rect 15616 19820 15650 19854
rect 15616 19752 15650 19786
rect 15616 19684 15650 19718
rect 15616 19616 15650 19650
rect 15616 19548 15650 19582
rect 15616 19480 15650 19514
rect 15616 19412 15650 19446
rect 15616 19344 15650 19378
rect 15616 19276 15650 19310
rect 15616 19208 15650 19242
rect 15616 19140 15650 19174
rect 14716 19020 14750 19106
rect 15616 19020 15650 19106
rect 14716 18986 14826 19020
rect 14860 18986 14894 19020
rect 14928 18986 14962 19020
rect 14996 18986 15030 19020
rect 15064 18986 15098 19020
rect 15132 18986 15166 19020
rect 15200 18986 15234 19020
rect 15268 18986 15302 19020
rect 15336 18986 15370 19020
rect 15404 18986 15438 19020
rect 15472 18986 15506 19020
rect 15540 18986 15650 19020
rect 15876 20100 15998 20134
rect 16032 20100 16066 20134
rect 16100 20100 16134 20134
rect 16168 20100 16202 20134
rect 16236 20100 16270 20134
rect 16304 20100 16426 20134
rect 15876 20019 15910 20100
rect 15876 19951 15910 19985
rect 16392 20019 16426 20100
rect 15876 19883 15910 19917
rect 15876 19815 15910 19849
rect 15876 19747 15910 19781
rect 15876 19679 15910 19713
rect 15876 19611 15910 19645
rect 15876 19543 15910 19577
rect 15876 19475 15910 19509
rect 15876 19407 15910 19441
rect 15876 19339 15910 19373
rect 15876 19271 15910 19305
rect 15876 19203 15910 19237
rect 15876 19135 15910 19169
rect 16392 19951 16426 19985
rect 16392 19883 16426 19917
rect 16392 19815 16426 19849
rect 16392 19747 16426 19781
rect 16392 19679 16426 19713
rect 16392 19611 16426 19645
rect 16392 19543 16426 19577
rect 16392 19475 16426 19509
rect 16392 19407 16426 19441
rect 16392 19339 16426 19373
rect 16392 19271 16426 19305
rect 16392 19203 16426 19237
rect 15876 19020 15910 19101
rect 16392 19135 16426 19169
rect 16392 19020 16426 19101
rect 15876 18986 15998 19020
rect 16032 18986 16066 19020
rect 16100 18986 16134 19020
rect 16168 18986 16202 19020
rect 16236 18986 16270 19020
rect 16304 18986 16426 19020
rect 16656 20067 16690 20101
rect 16656 19999 16690 20033
rect 16656 19931 16690 19965
rect 16656 19863 16690 19897
rect 16656 19795 16690 19829
rect 16656 19727 16690 19761
rect 16656 19659 16690 19693
rect 16656 19591 16690 19625
rect 16656 19523 16690 19557
rect 16656 19455 16690 19489
rect 16656 19387 16690 19421
rect 16656 19319 16690 19353
rect 16656 19251 16690 19285
rect 16656 19183 16690 19217
rect 16656 19115 16690 19149
rect 16656 19047 16690 19081
rect 13182 18871 13216 18905
rect 13182 18803 13216 18837
rect 14410 18939 14444 18973
rect 14410 18871 14444 18905
rect 13182 18735 13216 18769
rect 13182 18667 13216 18701
rect 13182 18599 13216 18633
rect 14410 18803 14444 18837
rect 14410 18735 14444 18769
rect 16656 18979 16690 19013
rect 16656 18911 16690 18945
rect 16952 21291 16986 21325
rect 16952 21223 16986 21257
rect 16952 21155 16986 21189
rect 16952 21087 16986 21121
rect 16952 21019 16986 21053
rect 16952 20951 16986 20985
rect 16952 20883 16986 20917
rect 16952 20815 16986 20849
rect 16952 20747 16986 20781
rect 16952 20679 16986 20713
rect 16952 20611 16986 20645
rect 16952 20543 16986 20577
rect 16952 20475 16986 20509
rect 16952 20407 16986 20441
rect 16952 20339 16986 20373
rect 16952 20271 16986 20305
rect 16952 20203 16986 20237
rect 16952 20135 16986 20169
rect 16952 20067 16986 20101
rect 16952 19999 16986 20033
rect 16952 19931 16986 19965
rect 16952 19863 16986 19897
rect 16952 19795 16986 19829
rect 16952 19727 16986 19761
rect 16952 19659 16986 19693
rect 16952 19591 16986 19625
rect 16952 19523 16986 19557
rect 16952 19455 16986 19489
rect 16952 19387 16986 19421
rect 16952 19319 16986 19353
rect 16952 19251 16986 19285
rect 16952 19183 16986 19217
rect 16952 19115 16986 19149
rect 16952 19047 16986 19081
rect 16952 18979 16986 19013
rect 16952 18911 16986 18945
rect 16656 18790 16690 18877
rect 16952 18790 16986 18877
rect 16656 18756 16770 18790
rect 16804 18756 16838 18790
rect 16872 18756 16986 18790
rect 17266 21466 17380 21500
rect 17414 21466 17448 21500
rect 17482 21466 17596 21500
rect 17266 21393 17300 21466
rect 17562 21393 17596 21466
rect 17266 21325 17300 21359
rect 17266 21257 17300 21291
rect 17266 21189 17300 21223
rect 17266 21121 17300 21155
rect 17266 21053 17300 21087
rect 17266 20985 17300 21019
rect 17266 20917 17300 20951
rect 17266 20849 17300 20883
rect 17266 20781 17300 20815
rect 17266 20713 17300 20747
rect 17266 20645 17300 20679
rect 17266 20577 17300 20611
rect 17266 20509 17300 20543
rect 17266 20441 17300 20475
rect 17266 20373 17300 20407
rect 17266 20305 17300 20339
rect 17266 20237 17300 20271
rect 17266 20169 17300 20203
rect 17266 20101 17300 20135
rect 17266 20033 17300 20067
rect 17266 19965 17300 19999
rect 17266 19897 17300 19931
rect 17266 19829 17300 19863
rect 17266 19761 17300 19795
rect 17266 19693 17300 19727
rect 17266 19625 17300 19659
rect 17266 19557 17300 19591
rect 17266 19489 17300 19523
rect 17266 19421 17300 19455
rect 17266 19353 17300 19387
rect 17266 19285 17300 19319
rect 17266 19217 17300 19251
rect 17266 19149 17300 19183
rect 17266 19081 17300 19115
rect 17266 19013 17300 19047
rect 17266 18945 17300 18979
rect 17266 18877 17300 18911
rect 17266 18809 17300 18843
rect 14410 18667 14444 18701
rect 17266 18741 17300 18775
rect 14410 18599 14444 18633
rect 13182 18531 13216 18565
rect 13182 18463 13216 18497
rect 14410 18531 14444 18565
rect 14410 18463 14444 18497
rect 13182 18395 13216 18429
rect 13182 18327 13216 18361
rect 13182 18259 13216 18293
rect 13182 18191 13216 18225
rect 14410 18395 14444 18429
rect 14410 18327 14444 18361
rect 14410 18259 14444 18293
rect 14410 18191 14444 18225
rect 13182 18123 13216 18157
rect 13182 18055 13216 18089
rect 14410 18123 14444 18157
rect 14410 18055 14444 18089
rect 13182 17987 13216 18021
rect 13182 17919 13216 17953
rect 13182 17851 13216 17885
rect 13182 17783 13216 17817
rect 14410 17987 14444 18021
rect 14902 18634 15026 18668
rect 15060 18634 15094 18668
rect 15128 18634 15252 18668
rect 14902 18547 14936 18634
rect 15218 18547 15252 18634
rect 14902 18479 14936 18513
rect 14902 18411 14936 18445
rect 14902 18343 14936 18377
rect 14902 18275 14936 18309
rect 14902 18207 14936 18241
rect 14902 18139 14936 18173
rect 14902 18071 14936 18105
rect 14902 18003 14936 18037
rect 14410 17919 14444 17953
rect 14410 17851 14444 17885
rect 13182 17715 13216 17749
rect 13182 17647 13216 17681
rect 14410 17783 14444 17817
rect 14410 17715 14444 17749
rect 13182 17579 13216 17613
rect 13182 17511 13216 17545
rect 13182 17443 13216 17477
rect 14410 17647 14444 17681
rect 14410 17579 14444 17613
rect 14410 17511 14444 17545
rect 14410 17443 14444 17477
rect 13182 17375 13216 17409
rect 13182 17307 13216 17341
rect 14410 17375 14444 17409
rect 14410 17307 14444 17341
rect 13182 17239 13216 17273
rect 13182 17171 13216 17205
rect 13182 17103 13216 17137
rect 13182 17035 13216 17069
rect 14410 17239 14444 17273
rect 14410 17171 14444 17205
rect 14410 17103 14444 17137
rect 14410 17035 14444 17069
rect 13182 16967 13216 17001
rect 13182 16899 13216 16933
rect 14410 16967 14444 17001
rect 14410 16899 14444 16933
rect 13182 16794 13216 16865
rect 14410 16794 14444 16865
rect 13182 16760 13286 16794
rect 13320 16760 13354 16794
rect 13388 16760 13422 16794
rect 13456 16760 13490 16794
rect 13524 16760 13558 16794
rect 13592 16760 13626 16794
rect 13660 16760 13694 16794
rect 13728 16760 13762 16794
rect 13796 16760 13830 16794
rect 13864 16760 13898 16794
rect 13932 16760 13966 16794
rect 14000 16760 14034 16794
rect 14068 16760 14102 16794
rect 14136 16760 14170 16794
rect 14204 16760 14238 16794
rect 14272 16760 14306 16794
rect 14340 16760 14444 16794
rect 14512 17950 14626 17984
rect 14660 17950 14694 17984
rect 14728 17950 14842 17984
rect 14512 17865 14546 17950
rect 14808 17865 14842 17950
rect 14512 17797 14546 17831
rect 14512 17729 14546 17763
rect 14512 17661 14546 17695
rect 14512 17593 14546 17627
rect 14512 17525 14546 17559
rect 14512 17457 14546 17491
rect 14512 17389 14546 17423
rect 14512 17321 14546 17355
rect 14512 17253 14546 17287
rect 14512 17185 14546 17219
rect 14512 17117 14546 17151
rect 14512 17049 14546 17083
rect 14512 16981 14546 17015
rect 14512 16913 14546 16947
rect 14808 17797 14842 17831
rect 14808 17729 14842 17763
rect 14808 17661 14842 17695
rect 14808 17593 14842 17627
rect 14808 17525 14842 17559
rect 14808 17457 14842 17491
rect 14808 17389 14842 17423
rect 14808 17321 14842 17355
rect 14808 17253 14842 17287
rect 14808 17185 14842 17219
rect 14808 17117 14842 17151
rect 14808 17049 14842 17083
rect 14808 16981 14842 17015
rect 14808 16913 14842 16947
rect 14512 16794 14546 16879
rect 14808 16794 14842 16879
rect 14512 16760 14626 16794
rect 14660 16760 14694 16794
rect 14728 16760 14842 16794
rect 14902 17935 14936 17969
rect 14902 17867 14936 17901
rect 14902 17799 14936 17833
rect 14902 17731 14936 17765
rect 14902 17663 14936 17697
rect 14902 17595 14936 17629
rect 14902 17527 14936 17561
rect 14902 17459 14936 17493
rect 14902 17391 14936 17425
rect 14902 17323 14936 17357
rect 14902 17255 14936 17289
rect 14902 17187 14936 17221
rect 14902 17119 14936 17153
rect 14902 17051 14936 17085
rect 14902 16983 14936 17017
rect 14902 16915 14936 16949
rect 15218 18479 15252 18513
rect 15218 18411 15252 18445
rect 15218 18343 15252 18377
rect 15218 18275 15252 18309
rect 15218 18207 15252 18241
rect 15218 18139 15252 18173
rect 15218 18071 15252 18105
rect 15218 18003 15252 18037
rect 15218 17935 15252 17969
rect 15218 17867 15252 17901
rect 15218 17799 15252 17833
rect 15218 17731 15252 17765
rect 15218 17663 15252 17697
rect 15218 17595 15252 17629
rect 15218 17527 15252 17561
rect 15218 17459 15252 17493
rect 15218 17391 15252 17425
rect 15218 17323 15252 17357
rect 15218 17255 15252 17289
rect 15218 17187 15252 17221
rect 15218 17119 15252 17153
rect 15218 17051 15252 17085
rect 15218 16983 15252 17017
rect 15218 16915 15252 16949
rect 14902 16794 14936 16881
rect 15218 16794 15252 16881
rect 14902 16760 15026 16794
rect 15060 16760 15094 16794
rect 15128 16760 15252 16794
rect 15312 18634 15436 18668
rect 15470 18634 15504 18668
rect 15538 18634 15662 18668
rect 15312 18547 15346 18634
rect 15628 18547 15662 18634
rect 15312 18479 15346 18513
rect 15312 18411 15346 18445
rect 15312 18343 15346 18377
rect 15312 18275 15346 18309
rect 15312 18207 15346 18241
rect 15312 18139 15346 18173
rect 15312 18071 15346 18105
rect 15312 18003 15346 18037
rect 15312 17935 15346 17969
rect 15312 17867 15346 17901
rect 15312 17799 15346 17833
rect 15312 17731 15346 17765
rect 15312 17663 15346 17697
rect 15312 17595 15346 17629
rect 15312 17527 15346 17561
rect 15312 17459 15346 17493
rect 15312 17391 15346 17425
rect 15312 17323 15346 17357
rect 15312 17255 15346 17289
rect 15312 17187 15346 17221
rect 15312 17119 15346 17153
rect 15312 17051 15346 17085
rect 15312 16983 15346 17017
rect 15312 16915 15346 16949
rect 15628 18479 15662 18513
rect 15628 18411 15662 18445
rect 15628 18343 15662 18377
rect 15628 18275 15662 18309
rect 15628 18207 15662 18241
rect 15628 18139 15662 18173
rect 15628 18071 15662 18105
rect 15628 18003 15662 18037
rect 16124 18651 16238 18685
rect 16272 18651 16306 18685
rect 16340 18651 16454 18685
rect 16124 18556 16158 18651
rect 16420 18556 16454 18651
rect 16124 18488 16158 18522
rect 16124 18420 16158 18454
rect 16124 18352 16158 18386
rect 16124 18284 16158 18318
rect 16124 18216 16158 18250
rect 16124 18148 16158 18182
rect 16124 18080 16158 18114
rect 16124 18012 16158 18046
rect 15628 17935 15662 17969
rect 15628 17867 15662 17901
rect 15628 17799 15662 17833
rect 15628 17731 15662 17765
rect 15628 17663 15662 17697
rect 15628 17595 15662 17629
rect 15628 17527 15662 17561
rect 15628 17459 15662 17493
rect 15628 17391 15662 17425
rect 15628 17323 15662 17357
rect 15628 17255 15662 17289
rect 15628 17187 15662 17221
rect 15628 17119 15662 17153
rect 15628 17051 15662 17085
rect 15628 16983 15662 17017
rect 15628 16915 15662 16949
rect 15312 16794 15346 16881
rect 15628 16794 15662 16881
rect 15312 16760 15436 16794
rect 15470 16760 15504 16794
rect 15538 16760 15662 16794
rect 15732 17950 15846 17984
rect 15880 17950 15914 17984
rect 15948 17950 16062 17984
rect 15732 17865 15766 17950
rect 16028 17865 16062 17950
rect 15732 17797 15766 17831
rect 15732 17729 15766 17763
rect 15732 17661 15766 17695
rect 15732 17593 15766 17627
rect 15732 17525 15766 17559
rect 15732 17457 15766 17491
rect 15732 17389 15766 17423
rect 15732 17321 15766 17355
rect 15732 17253 15766 17287
rect 15732 17185 15766 17219
rect 15732 17117 15766 17151
rect 15732 17049 15766 17083
rect 15732 16981 15766 17015
rect 15732 16913 15766 16947
rect 16028 17797 16062 17831
rect 16028 17729 16062 17763
rect 16028 17661 16062 17695
rect 16028 17593 16062 17627
rect 16028 17525 16062 17559
rect 16028 17457 16062 17491
rect 16028 17389 16062 17423
rect 16028 17321 16062 17355
rect 16028 17253 16062 17287
rect 16028 17185 16062 17219
rect 16028 17117 16062 17151
rect 16028 17049 16062 17083
rect 16028 16981 16062 17015
rect 16028 16913 16062 16947
rect 15732 16794 15766 16879
rect 16028 16794 16062 16879
rect 15732 16760 15846 16794
rect 15880 16760 15914 16794
rect 15948 16760 16062 16794
rect 16124 17944 16158 17978
rect 16124 17876 16158 17910
rect 16124 17808 16158 17842
rect 16124 17740 16158 17774
rect 16124 17672 16158 17706
rect 16124 17604 16158 17638
rect 16124 17536 16158 17570
rect 16124 17468 16158 17502
rect 16124 17400 16158 17434
rect 16124 17332 16158 17366
rect 16124 17264 16158 17298
rect 16124 17196 16158 17230
rect 16124 17128 16158 17162
rect 16124 17060 16158 17094
rect 16124 16992 16158 17026
rect 16124 16924 16158 16958
rect 16420 18488 16454 18522
rect 17266 18673 17300 18707
rect 17266 18605 17300 18639
rect 17266 18537 17300 18571
rect 17266 18469 17300 18503
rect 16420 18420 16454 18454
rect 16420 18352 16454 18386
rect 16420 18284 16454 18318
rect 16420 18216 16454 18250
rect 16420 18148 16454 18182
rect 16686 18426 16782 18460
rect 16816 18426 16850 18460
rect 16884 18426 16980 18460
rect 16686 18364 16720 18426
rect 16946 18364 16980 18426
rect 16686 18296 16720 18330
rect 16946 18296 16980 18330
rect 16686 18200 16720 18262
rect 16946 18200 16980 18262
rect 16686 18166 16782 18200
rect 16816 18166 16850 18200
rect 16884 18166 16980 18200
rect 17266 18401 17300 18435
rect 17266 18333 17300 18367
rect 17266 18265 17300 18299
rect 17266 18197 17300 18231
rect 16420 18080 16454 18114
rect 16420 18012 16454 18046
rect 16420 17944 16454 17978
rect 16420 17876 16454 17910
rect 16420 17808 16454 17842
rect 16420 17740 16454 17774
rect 16420 17672 16454 17706
rect 16420 17604 16454 17638
rect 16420 17536 16454 17570
rect 16420 17468 16454 17502
rect 16420 17400 16454 17434
rect 17266 18129 17300 18163
rect 17266 18061 17300 18095
rect 17266 17993 17300 18027
rect 17266 17925 17300 17959
rect 17266 17857 17300 17891
rect 17266 17789 17300 17823
rect 17266 17721 17300 17755
rect 17266 17653 17300 17687
rect 17266 17585 17300 17619
rect 17266 17517 17300 17551
rect 17562 21325 17596 21359
rect 17562 21257 17596 21291
rect 17562 21189 17596 21223
rect 17562 21121 17596 21155
rect 17562 21053 17596 21087
rect 17562 20985 17596 21019
rect 17562 20917 17596 20951
rect 17562 20849 17596 20883
rect 17562 20781 17596 20815
rect 17562 20713 17596 20747
rect 17562 20645 17596 20679
rect 17562 20577 17596 20611
rect 17562 20509 17596 20543
rect 17562 20441 17596 20475
rect 17562 20373 17596 20407
rect 17562 20305 17596 20339
rect 17562 20237 17596 20271
rect 17562 20169 17596 20203
rect 17562 20101 17596 20135
rect 17562 20033 17596 20067
rect 17562 19965 17596 19999
rect 17562 19897 17596 19931
rect 17562 19829 17596 19863
rect 17562 19761 17596 19795
rect 17562 19693 17596 19727
rect 17562 19625 17596 19659
rect 17562 19557 17596 19591
rect 17562 19489 17596 19523
rect 17562 19421 17596 19455
rect 17562 19353 17596 19387
rect 17562 19285 17596 19319
rect 17562 19217 17596 19251
rect 17562 19149 17596 19183
rect 17562 19081 17596 19115
rect 17562 19013 17596 19047
rect 17562 18945 17596 18979
rect 17562 18877 17596 18911
rect 17562 18809 17596 18843
rect 17562 18741 17596 18775
rect 17562 18673 17596 18707
rect 17562 18605 17596 18639
rect 17562 18537 17596 18571
rect 17562 18469 17596 18503
rect 17562 18401 17596 18435
rect 17562 18333 17596 18367
rect 17562 18265 17596 18299
rect 17562 18197 17596 18231
rect 17562 18129 17596 18163
rect 17562 18061 17596 18095
rect 17562 17993 17596 18027
rect 17562 17925 17596 17959
rect 17562 17857 17596 17891
rect 17562 17789 17596 17823
rect 17562 17721 17596 17755
rect 17562 17653 17596 17687
rect 17562 17585 17596 17619
rect 17562 17517 17596 17551
rect 17266 17410 17300 17483
rect 17562 17410 17596 17483
rect 17266 17376 17380 17410
rect 17414 17376 17448 17410
rect 17482 17376 17596 17410
rect 16420 17332 16454 17366
rect 16420 17264 16454 17298
rect 16420 17196 16454 17230
rect 16420 17128 16454 17162
rect 16420 17060 16454 17094
rect 16420 16992 16454 17026
rect 16420 16924 16454 16958
rect 16124 16795 16158 16890
rect 16420 16795 16454 16890
rect 16124 16761 16238 16795
rect 16272 16761 16306 16795
rect 16340 16761 16454 16795
rect 14308 16044 14432 16078
rect 14466 16044 14500 16078
rect 14534 16044 14568 16078
rect 14602 16044 14636 16078
rect 14670 16044 14704 16078
rect 14738 16044 14772 16078
rect 14806 16044 14840 16078
rect 14874 16044 14908 16078
rect 14942 16044 14976 16078
rect 15010 16044 15044 16078
rect 15078 16044 15112 16078
rect 15146 16044 15180 16078
rect 15214 16044 15338 16078
rect 14308 15975 14342 16044
rect 14308 15907 14342 15941
rect 15304 15975 15338 16044
rect 15304 15907 15338 15941
rect 14308 15839 14342 15873
rect 14308 15771 14342 15805
rect 14308 15703 14342 15737
rect 13458 15604 13582 15638
rect 13616 15604 13650 15638
rect 13684 15604 13808 15638
rect 13458 15517 13492 15604
rect 13774 15517 13808 15604
rect 13458 15449 13492 15483
rect 13458 15381 13492 15415
rect 13458 15313 13492 15347
rect 13458 15245 13492 15279
rect 13458 15177 13492 15211
rect 13458 15109 13492 15143
rect 13458 15041 13492 15075
rect 13458 14973 13492 15007
rect 13458 14905 13492 14939
rect 13458 14837 13492 14871
rect 13458 14769 13492 14803
rect 13458 14701 13492 14735
rect 13458 14633 13492 14667
rect 13458 14565 13492 14599
rect 13458 14497 13492 14531
rect 13458 14429 13492 14463
rect 13458 14361 13492 14395
rect 13458 14293 13492 14327
rect 13458 14225 13492 14259
rect 13458 14157 13492 14191
rect 13458 14089 13492 14123
rect 13458 14021 13492 14055
rect 13458 13953 13492 13987
rect 13458 13885 13492 13919
rect 13774 15449 13808 15483
rect 13774 15381 13808 15415
rect 13774 15313 13808 15347
rect 13774 15245 13808 15279
rect 13774 15177 13808 15211
rect 13774 15109 13808 15143
rect 13774 15041 13808 15075
rect 13774 14973 13808 15007
rect 13774 14905 13808 14939
rect 13774 14837 13808 14871
rect 13774 14769 13808 14803
rect 13774 14701 13808 14735
rect 13774 14633 13808 14667
rect 13774 14565 13808 14599
rect 13774 14497 13808 14531
rect 13774 14429 13808 14463
rect 13774 14361 13808 14395
rect 13774 14293 13808 14327
rect 13774 14225 13808 14259
rect 13774 14157 13808 14191
rect 13774 14089 13808 14123
rect 13774 14021 13808 14055
rect 13774 13953 13808 13987
rect 13774 13885 13808 13919
rect 13458 13764 13492 13851
rect 13774 13764 13808 13851
rect 13458 13730 13582 13764
rect 13616 13730 13650 13764
rect 13684 13730 13808 13764
rect 14308 15635 14342 15669
rect 14308 15567 14342 15601
rect 14308 15499 14342 15533
rect 14308 15431 14342 15465
rect 14308 15363 14342 15397
rect 14308 15295 14342 15329
rect 14308 15227 14342 15261
rect 14308 15159 14342 15193
rect 14308 15091 14342 15125
rect 14308 15023 14342 15057
rect 14308 14955 14342 14989
rect 14308 14887 14342 14921
rect 14308 14819 14342 14853
rect 14308 14751 14342 14785
rect 14308 14683 14342 14717
rect 14308 14615 14342 14649
rect 14308 14547 14342 14581
rect 14308 14479 14342 14513
rect 14308 14411 14342 14445
rect 14308 14343 14342 14377
rect 14308 14275 14342 14309
rect 14308 14207 14342 14241
rect 14308 14139 14342 14173
rect 14308 14071 14342 14105
rect 14308 14003 14342 14037
rect 14308 13935 14342 13969
rect 15304 15839 15338 15873
rect 15304 15771 15338 15805
rect 15304 15703 15338 15737
rect 15304 15635 15338 15669
rect 15304 15567 15338 15601
rect 15304 15499 15338 15533
rect 15304 15431 15338 15465
rect 15304 15363 15338 15397
rect 15304 15295 15338 15329
rect 15304 15227 15338 15261
rect 15304 15159 15338 15193
rect 15304 15091 15338 15125
rect 15304 15023 15338 15057
rect 15304 14955 15338 14989
rect 15304 14887 15338 14921
rect 15304 14819 15338 14853
rect 15304 14751 15338 14785
rect 15304 14683 15338 14717
rect 15304 14615 15338 14649
rect 15304 14547 15338 14581
rect 15304 14479 15338 14513
rect 15304 14411 15338 14445
rect 15304 14343 15338 14377
rect 15304 14275 15338 14309
rect 15304 14207 15338 14241
rect 15304 14139 15338 14173
rect 15304 14071 15338 14105
rect 15304 14003 15338 14037
rect 15304 13935 15338 13969
rect 14308 13867 14342 13901
rect 14308 13764 14342 13833
rect 15304 13867 15338 13901
rect 15304 13764 15338 13833
rect 14308 13730 14432 13764
rect 14466 13730 14500 13764
rect 14534 13730 14568 13764
rect 14602 13730 14636 13764
rect 14670 13730 14704 13764
rect 14738 13730 14772 13764
rect 14806 13730 14840 13764
rect 14874 13730 14908 13764
rect 14942 13730 14976 13764
rect 15010 13730 15044 13764
rect 15078 13730 15112 13764
rect 15146 13730 15180 13764
rect 15214 13730 15338 13764
rect 16018 16060 16132 16094
rect 16166 16060 16200 16094
rect 16234 16060 16348 16094
rect 16018 15983 16052 16060
rect 16314 15983 16348 16060
rect 16018 15915 16052 15949
rect 16018 15847 16052 15881
rect 16018 15779 16052 15813
rect 16018 15711 16052 15745
rect 16018 15643 16052 15677
rect 16018 15575 16052 15609
rect 16018 15507 16052 15541
rect 16018 15439 16052 15473
rect 16018 15371 16052 15405
rect 16018 15303 16052 15337
rect 16018 15235 16052 15269
rect 16018 15167 16052 15201
rect 16018 15099 16052 15133
rect 16018 15031 16052 15065
rect 16018 14963 16052 14997
rect 16018 14895 16052 14929
rect 16018 14827 16052 14861
rect 16018 14759 16052 14793
rect 16018 14691 16052 14725
rect 16018 14623 16052 14657
rect 16018 14555 16052 14589
rect 16018 14487 16052 14521
rect 16018 14419 16052 14453
rect 16018 14351 16052 14385
rect 16018 14283 16052 14317
rect 16018 14215 16052 14249
rect 16018 14147 16052 14181
rect 16018 14079 16052 14113
rect 16018 14011 16052 14045
rect 16018 13943 16052 13977
rect 16018 13875 16052 13909
rect 16314 15915 16348 15949
rect 16314 15847 16348 15881
rect 16314 15779 16348 15813
rect 16314 15711 16348 15745
rect 16314 15643 16348 15677
rect 16314 15575 16348 15609
rect 16314 15507 16348 15541
rect 16314 15439 16348 15473
rect 16314 15371 16348 15405
rect 16314 15303 16348 15337
rect 16314 15235 16348 15269
rect 16314 15167 16348 15201
rect 16314 15099 16348 15133
rect 16314 15031 16348 15065
rect 16314 14963 16348 14997
rect 16314 14895 16348 14929
rect 16314 14827 16348 14861
rect 16314 14759 16348 14793
rect 16314 14691 16348 14725
rect 16314 14623 16348 14657
rect 16314 14555 16348 14589
rect 16314 14487 16348 14521
rect 16314 14419 16348 14453
rect 16314 14351 16348 14385
rect 16314 14283 16348 14317
rect 16314 14215 16348 14249
rect 16314 14147 16348 14181
rect 16314 14079 16348 14113
rect 16314 14011 16348 14045
rect 16314 13943 16348 13977
rect 16314 13875 16348 13909
rect 16018 13764 16052 13841
rect 16314 13764 16348 13841
rect 16018 13730 16132 13764
rect 16166 13730 16200 13764
rect 16234 13730 16348 13764
rect 13074 13546 17870 13590
rect 13074 13512 13329 13546
rect 13363 13512 13397 13546
rect 13431 13512 13465 13546
rect 13499 13512 13533 13546
rect 13567 13512 13601 13546
rect 13635 13512 13669 13546
rect 13703 13512 13737 13546
rect 13771 13512 13805 13546
rect 13839 13512 13873 13546
rect 13907 13512 13941 13546
rect 13975 13512 14009 13546
rect 14043 13512 14077 13546
rect 14111 13512 14145 13546
rect 14179 13512 14213 13546
rect 14247 13512 14281 13546
rect 14315 13512 14349 13546
rect 14383 13512 14417 13546
rect 14451 13512 14485 13546
rect 14519 13512 14553 13546
rect 14587 13512 14621 13546
rect 14655 13512 14689 13546
rect 14723 13512 14757 13546
rect 14791 13512 14825 13546
rect 14859 13512 14893 13546
rect 14927 13512 14961 13546
rect 14995 13512 15029 13546
rect 15063 13512 15097 13546
rect 15131 13512 15165 13546
rect 15199 13512 15233 13546
rect 15267 13512 15301 13546
rect 15335 13512 15369 13546
rect 15403 13512 15437 13546
rect 15471 13512 15505 13546
rect 15539 13512 15573 13546
rect 15607 13512 15641 13546
rect 15675 13512 15709 13546
rect 15743 13512 15777 13546
rect 15811 13512 15845 13546
rect 15879 13512 15913 13546
rect 15947 13512 15981 13546
rect 16015 13512 16049 13546
rect 16083 13512 16117 13546
rect 16151 13512 16185 13546
rect 16219 13512 16253 13546
rect 16287 13512 16321 13546
rect 16355 13512 16389 13546
rect 16423 13512 16457 13546
rect 16491 13512 16525 13546
rect 16559 13512 16593 13546
rect 16627 13512 16661 13546
rect 16695 13512 16729 13546
rect 16763 13512 16797 13546
rect 16831 13512 16865 13546
rect 16899 13512 16933 13546
rect 16967 13512 17001 13546
rect 17035 13512 17069 13546
rect 17103 13512 17137 13546
rect 17171 13512 17205 13546
rect 17239 13512 17273 13546
rect 17307 13512 17341 13546
rect 17375 13512 17409 13546
rect 17443 13512 17477 13546
rect 17511 13512 17545 13546
rect 17579 13512 17870 13546
rect 13074 13455 17870 13512
rect 13074 13416 13209 13455
rect 13074 13382 13122 13416
rect 13156 13382 13209 13416
rect 13074 13348 13209 13382
rect 13074 13314 13122 13348
rect 13156 13314 13209 13348
rect 17728 13425 17870 13455
rect 17728 13391 17785 13425
rect 17819 13391 17870 13425
rect 17728 13357 17870 13391
rect 13074 13280 13209 13314
rect 13074 13246 13122 13280
rect 13156 13246 13209 13280
rect 13074 13212 13209 13246
rect 13074 13178 13122 13212
rect 13156 13178 13209 13212
rect 13074 13144 13209 13178
rect 13074 13110 13122 13144
rect 13156 13110 13209 13144
rect 13074 13076 13209 13110
rect 13074 13042 13122 13076
rect 13156 13042 13209 13076
rect 17728 13323 17785 13357
rect 17819 13323 17870 13357
rect 17728 13289 17870 13323
rect 17728 13255 17785 13289
rect 17819 13255 17870 13289
rect 17728 13221 17870 13255
rect 17728 13187 17785 13221
rect 17819 13187 17870 13221
rect 17728 13153 17870 13187
rect 17728 13119 17785 13153
rect 17819 13119 17870 13153
rect 17728 13085 17870 13119
rect 13074 13008 13209 13042
rect 13074 12974 13122 13008
rect 13156 12974 13209 13008
rect 13074 12940 13209 12974
rect 13074 12906 13122 12940
rect 13156 12906 13209 12940
rect 13074 12872 13209 12906
rect 13074 12838 13122 12872
rect 13156 12838 13209 12872
rect 13074 12804 13209 12838
rect 13074 12770 13122 12804
rect 13156 12770 13209 12804
rect 13074 12736 13209 12770
rect 13074 12702 13122 12736
rect 13156 12702 13209 12736
rect 13074 12668 13209 12702
rect 13074 12634 13122 12668
rect 13156 12634 13209 12668
rect 13074 12600 13209 12634
rect 13074 12566 13122 12600
rect 13156 12566 13209 12600
rect 13074 12532 13209 12566
rect 13074 12498 13122 12532
rect 13156 12498 13209 12532
rect 13074 12464 13209 12498
rect 13074 12430 13122 12464
rect 13156 12430 13209 12464
rect 13074 12396 13209 12430
rect 13074 12362 13122 12396
rect 13156 12362 13209 12396
rect 13074 12328 13209 12362
rect 13074 12294 13122 12328
rect 13156 12294 13209 12328
rect 13074 12260 13209 12294
rect 13074 12226 13122 12260
rect 13156 12226 13209 12260
rect 13074 12192 13209 12226
rect 13074 12158 13122 12192
rect 13156 12158 13209 12192
rect 13074 12124 13209 12158
rect 13074 12090 13122 12124
rect 13156 12090 13209 12124
rect 13074 12056 13209 12090
rect 13074 12022 13122 12056
rect 13156 12022 13209 12056
rect 13074 11988 13209 12022
rect 13074 11954 13122 11988
rect 13156 11954 13209 11988
rect 13074 11920 13209 11954
rect 13074 11886 13122 11920
rect 13156 11886 13209 11920
rect 13074 11852 13209 11886
rect 13074 11818 13122 11852
rect 13156 11818 13209 11852
rect 13074 11784 13209 11818
rect 13074 11750 13122 11784
rect 13156 11750 13209 11784
rect 13074 11716 13209 11750
rect 13074 11682 13122 11716
rect 13156 11682 13209 11716
rect 13074 11648 13209 11682
rect 13074 11614 13122 11648
rect 13156 11614 13209 11648
rect 13074 11580 13209 11614
rect 13074 11546 13122 11580
rect 13156 11546 13209 11580
rect 13074 11512 13209 11546
rect 13074 11478 13122 11512
rect 13156 11478 13209 11512
rect 13074 11444 13209 11478
rect 13074 11410 13122 11444
rect 13156 11410 13209 11444
rect 13074 11376 13209 11410
rect 13074 11342 13122 11376
rect 13156 11342 13209 11376
rect 13074 11308 13209 11342
rect 13074 11274 13122 11308
rect 13156 11274 13209 11308
rect 13074 11240 13209 11274
rect 13074 11206 13122 11240
rect 13156 11206 13209 11240
rect 13074 11172 13209 11206
rect 13074 11138 13122 11172
rect 13156 11138 13209 11172
rect 13074 11104 13209 11138
rect 13074 11070 13122 11104
rect 13156 11070 13209 11104
rect 17728 13051 17785 13085
rect 17819 13051 17870 13085
rect 17728 13017 17870 13051
rect 17728 12983 17785 13017
rect 17819 12983 17870 13017
rect 17728 12949 17870 12983
rect 17728 12915 17785 12949
rect 17819 12915 17870 12949
rect 17728 12881 17870 12915
rect 17728 12847 17785 12881
rect 17819 12847 17870 12881
rect 17728 12813 17870 12847
rect 17728 12779 17785 12813
rect 17819 12779 17870 12813
rect 17728 12745 17870 12779
rect 17728 12711 17785 12745
rect 17819 12711 17870 12745
rect 17728 12677 17870 12711
rect 17728 12643 17785 12677
rect 17819 12643 17870 12677
rect 17728 12609 17870 12643
rect 17728 12575 17785 12609
rect 17819 12575 17870 12609
rect 17728 12541 17870 12575
rect 17728 12507 17785 12541
rect 17819 12507 17870 12541
rect 17728 12473 17870 12507
rect 17728 12439 17785 12473
rect 17819 12439 17870 12473
rect 17728 12405 17870 12439
rect 17728 12371 17785 12405
rect 17819 12371 17870 12405
rect 17728 12337 17870 12371
rect 17728 12303 17785 12337
rect 17819 12303 17870 12337
rect 17728 12269 17870 12303
rect 17728 12235 17785 12269
rect 17819 12235 17870 12269
rect 17728 12201 17870 12235
rect 17728 12167 17785 12201
rect 17819 12167 17870 12201
rect 17728 12133 17870 12167
rect 17728 12099 17785 12133
rect 17819 12099 17870 12133
rect 17728 12065 17870 12099
rect 17728 12031 17785 12065
rect 17819 12031 17870 12065
rect 17728 11997 17870 12031
rect 17728 11963 17785 11997
rect 17819 11963 17870 11997
rect 17728 11929 17870 11963
rect 17728 11895 17785 11929
rect 17819 11895 17870 11929
rect 17728 11861 17870 11895
rect 17728 11827 17785 11861
rect 17819 11827 17870 11861
rect 17728 11793 17870 11827
rect 17728 11759 17785 11793
rect 17819 11759 17870 11793
rect 17728 11725 17870 11759
rect 17728 11691 17785 11725
rect 17819 11691 17870 11725
rect 17728 11657 17870 11691
rect 17728 11623 17785 11657
rect 17819 11623 17870 11657
rect 17728 11589 17870 11623
rect 17728 11555 17785 11589
rect 17819 11555 17870 11589
rect 17728 11521 17870 11555
rect 17728 11487 17785 11521
rect 17819 11487 17870 11521
rect 17728 11453 17870 11487
rect 17728 11419 17785 11453
rect 17819 11419 17870 11453
rect 17728 11385 17870 11419
rect 17728 11351 17785 11385
rect 17819 11351 17870 11385
rect 17728 11317 17870 11351
rect 17728 11283 17785 11317
rect 17819 11283 17870 11317
rect 17728 11249 17870 11283
rect 17728 11215 17785 11249
rect 17819 11215 17870 11249
rect 17728 11181 17870 11215
rect 17728 11147 17785 11181
rect 17819 11147 17870 11181
rect 17728 11113 17870 11147
rect 17728 11079 17785 11113
rect 17819 11079 17870 11113
rect 13074 11036 13209 11070
rect 13074 11002 13122 11036
rect 13156 11002 13209 11036
rect 13074 10968 13209 11002
rect 13074 10934 13122 10968
rect 13156 10934 13209 10968
rect 13074 10900 13209 10934
rect 17728 11045 17870 11079
rect 13074 10866 13122 10900
rect 13156 10866 13209 10900
rect 17728 11011 17785 11045
rect 17819 11011 17870 11045
rect 17728 10977 17870 11011
rect 17728 10943 17785 10977
rect 17819 10943 17870 10977
rect 17728 10909 17870 10943
rect 13074 10832 13209 10866
rect 13074 10798 13122 10832
rect 13156 10798 13209 10832
rect 13074 10738 13209 10798
rect 17728 10875 17785 10909
rect 17819 10875 17870 10909
rect 17728 10841 17870 10875
rect 17728 10807 17785 10841
rect 17819 10807 17870 10841
rect 17728 10738 17870 10807
rect 13074 10693 17870 10738
rect 13074 10659 13371 10693
rect 13405 10659 13439 10693
rect 13473 10659 13507 10693
rect 13541 10659 13575 10693
rect 13609 10659 13643 10693
rect 13677 10659 13711 10693
rect 13745 10659 13779 10693
rect 13813 10659 13847 10693
rect 13881 10659 13915 10693
rect 13949 10659 13983 10693
rect 14017 10659 14051 10693
rect 14085 10659 14119 10693
rect 14153 10659 14187 10693
rect 14221 10659 14255 10693
rect 14289 10659 14323 10693
rect 14357 10659 14391 10693
rect 14425 10659 14459 10693
rect 14493 10659 14527 10693
rect 14561 10659 14595 10693
rect 14629 10659 14663 10693
rect 14697 10659 14731 10693
rect 14765 10659 14799 10693
rect 14833 10659 14867 10693
rect 14901 10659 14935 10693
rect 14969 10659 15003 10693
rect 15037 10659 15071 10693
rect 15105 10659 15139 10693
rect 15173 10659 15207 10693
rect 15241 10659 15275 10693
rect 15309 10659 15343 10693
rect 15377 10659 15411 10693
rect 15445 10659 15479 10693
rect 15513 10659 15547 10693
rect 15581 10659 15615 10693
rect 15649 10659 15683 10693
rect 15717 10659 15751 10693
rect 15785 10659 15819 10693
rect 15853 10659 15887 10693
rect 15921 10659 15955 10693
rect 15989 10659 16023 10693
rect 16057 10659 16091 10693
rect 16125 10659 16159 10693
rect 16193 10659 16227 10693
rect 16261 10659 16295 10693
rect 16329 10659 16363 10693
rect 16397 10659 16431 10693
rect 16465 10659 16499 10693
rect 16533 10659 16567 10693
rect 16601 10659 16635 10693
rect 16669 10659 16703 10693
rect 16737 10659 16771 10693
rect 16805 10659 16839 10693
rect 16873 10659 16907 10693
rect 16941 10659 16975 10693
rect 17009 10659 17043 10693
rect 17077 10659 17111 10693
rect 17145 10659 17179 10693
rect 17213 10659 17247 10693
rect 17281 10659 17315 10693
rect 17349 10659 17383 10693
rect 17417 10659 17451 10693
rect 17485 10659 17519 10693
rect 17553 10659 17587 10693
rect 17621 10659 17870 10693
rect 13074 10610 17870 10659
<< nsubdiff >>
rect 15716 23338 15838 23372
rect 15872 23338 15906 23372
rect 15940 23338 15974 23372
rect 16008 23338 16042 23372
rect 16076 23338 16110 23372
rect 16144 23338 16266 23372
rect 15716 23260 15750 23338
rect 15716 23192 15750 23226
rect 16232 23260 16266 23338
rect 16232 23192 16266 23226
rect 15716 23124 15750 23158
rect 15716 23056 15750 23090
rect 15716 22988 15750 23022
rect 15716 22920 15750 22954
rect 15716 22852 15750 22886
rect 15716 22784 15750 22818
rect 15716 22716 15750 22750
rect 15716 22648 15750 22682
rect 15716 22580 15750 22614
rect 15716 22512 15750 22546
rect 15716 22444 15750 22478
rect 15716 22376 15750 22410
rect 15716 22308 15750 22342
rect 15716 22240 15750 22274
rect 15716 22172 15750 22206
rect 15716 22104 15750 22138
rect 15716 22036 15750 22070
rect 15716 21968 15750 22002
rect 15716 21900 15750 21934
rect 15716 21832 15750 21866
rect 15716 21764 15750 21798
rect 15716 21696 15750 21730
rect 15716 21628 15750 21662
rect 15716 21560 15750 21594
rect 15716 21492 15750 21526
rect 15716 21424 15750 21458
rect 15716 21356 15750 21390
rect 15716 21288 15750 21322
rect 15716 21220 15750 21254
rect 16232 23124 16266 23158
rect 16232 23056 16266 23090
rect 16232 22988 16266 23022
rect 16232 22920 16266 22954
rect 16232 22852 16266 22886
rect 16232 22784 16266 22818
rect 16232 22716 16266 22750
rect 16232 22648 16266 22682
rect 16232 22580 16266 22614
rect 16232 22512 16266 22546
rect 16232 22444 16266 22478
rect 16232 22376 16266 22410
rect 16232 22308 16266 22342
rect 16232 22240 16266 22274
rect 16232 22172 16266 22206
rect 16232 22104 16266 22138
rect 16232 22036 16266 22070
rect 16232 21968 16266 22002
rect 16232 21900 16266 21934
rect 16232 21832 16266 21866
rect 16232 21764 16266 21798
rect 16232 21696 16266 21730
rect 16232 21628 16266 21662
rect 16232 21560 16266 21594
rect 16232 21492 16266 21526
rect 16232 21424 16266 21458
rect 16232 21356 16266 21390
rect 16232 21288 16266 21322
rect 16232 21220 16266 21254
rect 15716 21152 15750 21186
rect 15716 21040 15750 21118
rect 16232 21152 16266 21186
rect 16232 21040 16266 21118
rect 15716 21006 15838 21040
rect 15872 21006 15906 21040
rect 15940 21006 15974 21040
rect 16008 21006 16042 21040
rect 16076 21006 16110 21040
rect 16144 21006 16266 21040
rect 16978 16092 17100 16126
rect 17134 16092 17168 16126
rect 17202 16092 17236 16126
rect 17270 16092 17304 16126
rect 17338 16092 17372 16126
rect 17406 16092 17528 16126
rect 16978 16014 17012 16092
rect 16978 15946 17012 15980
rect 17494 16014 17528 16092
rect 17494 15946 17528 15980
rect 16978 15878 17012 15912
rect 16978 15810 17012 15844
rect 16978 15742 17012 15776
rect 16978 15674 17012 15708
rect 16978 15606 17012 15640
rect 16978 15538 17012 15572
rect 16978 15470 17012 15504
rect 16978 15402 17012 15436
rect 16978 15334 17012 15368
rect 16978 15266 17012 15300
rect 16978 15198 17012 15232
rect 16978 15130 17012 15164
rect 16978 15062 17012 15096
rect 16978 14994 17012 15028
rect 16978 14926 17012 14960
rect 16978 14858 17012 14892
rect 16978 14790 17012 14824
rect 16978 14722 17012 14756
rect 16978 14654 17012 14688
rect 16978 14586 17012 14620
rect 16978 14518 17012 14552
rect 16978 14450 17012 14484
rect 16978 14382 17012 14416
rect 16978 14314 17012 14348
rect 16978 14246 17012 14280
rect 16978 14178 17012 14212
rect 16978 14110 17012 14144
rect 16978 14042 17012 14076
rect 16978 13974 17012 14008
rect 17494 15878 17528 15912
rect 17494 15810 17528 15844
rect 17494 15742 17528 15776
rect 17494 15674 17528 15708
rect 17494 15606 17528 15640
rect 17494 15538 17528 15572
rect 17494 15470 17528 15504
rect 17494 15402 17528 15436
rect 17494 15334 17528 15368
rect 17494 15266 17528 15300
rect 17494 15198 17528 15232
rect 17494 15130 17528 15164
rect 17494 15062 17528 15096
rect 17494 14994 17528 15028
rect 17494 14926 17528 14960
rect 17494 14858 17528 14892
rect 17494 14790 17528 14824
rect 17494 14722 17528 14756
rect 17494 14654 17528 14688
rect 17494 14586 17528 14620
rect 17494 14518 17528 14552
rect 17494 14450 17528 14484
rect 17494 14382 17528 14416
rect 17494 14314 17528 14348
rect 17494 14246 17528 14280
rect 17494 14178 17528 14212
rect 17494 14110 17528 14144
rect 17494 14042 17528 14076
rect 17494 13974 17528 14008
rect 16978 13906 17012 13940
rect 16978 13794 17012 13872
rect 17494 13906 17528 13940
rect 17494 13794 17528 13872
rect 16978 13760 17100 13794
rect 17134 13760 17168 13794
rect 17202 13760 17236 13794
rect 17270 13760 17304 13794
rect 17338 13760 17372 13794
rect 17406 13760 17528 13794
<< psubdiffcont >>
rect 13023 24712 13057 24746
rect 13091 24712 13125 24746
rect 13159 24712 13193 24746
rect 13227 24712 13261 24746
rect 13295 24712 13329 24746
rect 13363 24712 13397 24746
rect 13431 24712 13465 24746
rect 13499 24712 13533 24746
rect 13567 24712 13601 24746
rect 13635 24712 13669 24746
rect 13703 24712 13737 24746
rect 13771 24712 13805 24746
rect 13839 24712 13873 24746
rect 13907 24712 13941 24746
rect 13975 24712 14009 24746
rect 14043 24712 14077 24746
rect 14111 24712 14145 24746
rect 14179 24712 14213 24746
rect 14247 24712 14281 24746
rect 14315 24712 14349 24746
rect 14383 24712 14417 24746
rect 14451 24712 14485 24746
rect 14519 24712 14553 24746
rect 14587 24712 14621 24746
rect 14655 24712 14689 24746
rect 14723 24712 14757 24746
rect 14791 24712 14825 24746
rect 14859 24712 14893 24746
rect 14927 24712 14961 24746
rect 14995 24712 15029 24746
rect 15063 24712 15097 24746
rect 15131 24712 15165 24746
rect 15199 24712 15233 24746
rect 15267 24712 15301 24746
rect 15335 24712 15369 24746
rect 15403 24712 15437 24746
rect 15471 24712 15505 24746
rect 15539 24712 15573 24746
rect 15607 24712 15641 24746
rect 15675 24712 15709 24746
rect 15743 24712 15777 24746
rect 15811 24712 15845 24746
rect 15879 24712 15913 24746
rect 15947 24712 15981 24746
rect 16015 24712 16049 24746
rect 16083 24712 16117 24746
rect 16151 24712 16185 24746
rect 16219 24712 16253 24746
rect 16287 24712 16321 24746
rect 16355 24712 16389 24746
rect 16423 24712 16457 24746
rect 16491 24712 16525 24746
rect 16559 24712 16593 24746
rect 16627 24712 16661 24746
rect 16695 24712 16729 24746
rect 16763 24712 16797 24746
rect 16831 24712 16865 24746
rect 16899 24712 16933 24746
rect 12916 24598 12950 24632
rect 12916 24530 12950 24564
rect 17006 24598 17040 24632
rect 17006 24530 17040 24564
rect 13023 24416 13057 24450
rect 13091 24416 13125 24450
rect 13159 24416 13193 24450
rect 13227 24416 13261 24450
rect 13295 24416 13329 24450
rect 13363 24416 13397 24450
rect 13431 24416 13465 24450
rect 13499 24416 13533 24450
rect 13567 24416 13601 24450
rect 13635 24416 13669 24450
rect 13703 24416 13737 24450
rect 13771 24416 13805 24450
rect 13839 24416 13873 24450
rect 13907 24416 13941 24450
rect 13975 24416 14009 24450
rect 14043 24416 14077 24450
rect 14111 24416 14145 24450
rect 14179 24416 14213 24450
rect 14247 24416 14281 24450
rect 14315 24416 14349 24450
rect 14383 24416 14417 24450
rect 14451 24416 14485 24450
rect 14519 24416 14553 24450
rect 14587 24416 14621 24450
rect 14655 24416 14689 24450
rect 14723 24416 14757 24450
rect 14791 24416 14825 24450
rect 14859 24416 14893 24450
rect 14927 24416 14961 24450
rect 14995 24416 15029 24450
rect 15063 24416 15097 24450
rect 15131 24416 15165 24450
rect 15199 24416 15233 24450
rect 15267 24416 15301 24450
rect 15335 24416 15369 24450
rect 15403 24416 15437 24450
rect 15471 24416 15505 24450
rect 15539 24416 15573 24450
rect 15607 24416 15641 24450
rect 15675 24416 15709 24450
rect 15743 24416 15777 24450
rect 15811 24416 15845 24450
rect 15879 24416 15913 24450
rect 15947 24416 15981 24450
rect 16015 24416 16049 24450
rect 16083 24416 16117 24450
rect 16151 24416 16185 24450
rect 16219 24416 16253 24450
rect 16287 24416 16321 24450
rect 16355 24416 16389 24450
rect 16423 24416 16457 24450
rect 16491 24416 16525 24450
rect 16559 24416 16593 24450
rect 16627 24416 16661 24450
rect 16695 24416 16729 24450
rect 16763 24416 16797 24450
rect 16831 24416 16865 24450
rect 16899 24416 16933 24450
rect 16666 24180 16700 24214
rect 16734 24180 16768 24214
rect 16802 24180 16836 24214
rect 16870 24180 16904 24214
rect 16938 24180 16972 24214
rect 17006 24180 17040 24214
rect 17074 24180 17108 24214
rect 17142 24180 17176 24214
rect 17210 24180 17244 24214
rect 17278 24180 17312 24214
rect 17346 24180 17380 24214
rect 17414 24180 17448 24214
rect 17482 24180 17516 24214
rect 17550 24180 17584 24214
rect 17618 24180 17652 24214
rect 16548 24077 16582 24111
rect 13075 24032 13109 24066
rect 13143 24032 13177 24066
rect 13211 24032 13245 24066
rect 13279 24032 13313 24066
rect 13347 24032 13381 24066
rect 13415 24032 13449 24066
rect 13483 24032 13517 24066
rect 13551 24032 13585 24066
rect 13619 24032 13653 24066
rect 13687 24032 13721 24066
rect 13755 24032 13789 24066
rect 13823 24032 13857 24066
rect 13891 24032 13925 24066
rect 13959 24032 13993 24066
rect 14027 24032 14061 24066
rect 14095 24032 14129 24066
rect 14163 24032 14197 24066
rect 14231 24032 14265 24066
rect 14299 24032 14333 24066
rect 14367 24032 14401 24066
rect 14435 24032 14469 24066
rect 14503 24032 14537 24066
rect 14571 24032 14605 24066
rect 14639 24032 14673 24066
rect 14707 24032 14741 24066
rect 12946 23918 12980 23952
rect 12946 23850 12980 23884
rect 14836 23918 14870 23952
rect 14836 23850 14870 23884
rect 13075 23736 13109 23770
rect 13143 23736 13177 23770
rect 13211 23736 13245 23770
rect 13279 23736 13313 23770
rect 13347 23736 13381 23770
rect 13415 23736 13449 23770
rect 13483 23736 13517 23770
rect 13551 23736 13585 23770
rect 13619 23736 13653 23770
rect 13687 23736 13721 23770
rect 13755 23736 13789 23770
rect 13823 23736 13857 23770
rect 13891 23736 13925 23770
rect 13959 23736 13993 23770
rect 14027 23736 14061 23770
rect 14095 23736 14129 23770
rect 14163 23736 14197 23770
rect 14231 23736 14265 23770
rect 14299 23736 14333 23770
rect 14367 23736 14401 23770
rect 14435 23736 14469 23770
rect 14503 23736 14537 23770
rect 14571 23736 14605 23770
rect 14639 23736 14673 23770
rect 14707 23736 14741 23770
rect 16548 24009 16582 24043
rect 17736 24077 17770 24111
rect 16548 23941 16582 23975
rect 16548 23873 16582 23907
rect 16548 23805 16582 23839
rect 16548 23737 16582 23771
rect 16548 23669 16582 23703
rect 16548 23601 16582 23635
rect 16548 23533 16582 23567
rect 16548 23465 16582 23499
rect 16548 23397 16582 23431
rect 15290 23326 15324 23360
rect 15358 23326 15392 23360
rect 13980 23290 14014 23324
rect 14048 23290 14082 23324
rect 14116 23290 14150 23324
rect 14184 23290 14218 23324
rect 14252 23290 14286 23324
rect 14320 23290 14354 23324
rect 14388 23290 14422 23324
rect 14456 23290 14490 23324
rect 14524 23290 14558 23324
rect 14592 23290 14626 23324
rect 14660 23290 14694 23324
rect 14728 23290 14762 23324
rect 13856 23187 13890 23221
rect 13856 23119 13890 23153
rect 14852 23187 14886 23221
rect 13856 23051 13890 23085
rect 13856 22983 13890 23017
rect 13856 22915 13890 22949
rect 13856 22847 13890 22881
rect 13856 22779 13890 22813
rect 13856 22711 13890 22745
rect 13856 22643 13890 22677
rect 13856 22575 13890 22609
rect 13856 22507 13890 22541
rect 13856 22439 13890 22473
rect 13856 22371 13890 22405
rect 13856 22303 13890 22337
rect 13856 22235 13890 22269
rect 13470 22166 13504 22200
rect 13538 22166 13572 22200
rect 13356 22047 13390 22081
rect 13356 21979 13390 22013
rect 13356 21911 13390 21945
rect 13356 21843 13390 21877
rect 13356 21775 13390 21809
rect 13356 21707 13390 21741
rect 13356 21639 13390 21673
rect 13356 21571 13390 21605
rect 13356 21503 13390 21537
rect 13356 21435 13390 21469
rect 13356 21367 13390 21401
rect 13356 21299 13390 21333
rect 13356 21231 13390 21265
rect 13356 21163 13390 21197
rect 13356 21095 13390 21129
rect 13652 22047 13686 22081
rect 13652 21979 13686 22013
rect 13652 21911 13686 21945
rect 13652 21843 13686 21877
rect 13652 21775 13686 21809
rect 13652 21707 13686 21741
rect 13652 21639 13686 21673
rect 13652 21571 13686 21605
rect 13652 21503 13686 21537
rect 13652 21435 13686 21469
rect 13652 21367 13686 21401
rect 13652 21299 13686 21333
rect 13652 21231 13686 21265
rect 13652 21163 13686 21197
rect 13652 21095 13686 21129
rect 13470 20976 13504 21010
rect 13538 20976 13572 21010
rect 13856 22167 13890 22201
rect 13856 22099 13890 22133
rect 13856 22031 13890 22065
rect 13856 21963 13890 21997
rect 13856 21895 13890 21929
rect 13856 21827 13890 21861
rect 13856 21759 13890 21793
rect 13856 21691 13890 21725
rect 13856 21623 13890 21657
rect 13856 21555 13890 21589
rect 13856 21487 13890 21521
rect 13856 21419 13890 21453
rect 13856 21351 13890 21385
rect 13856 21283 13890 21317
rect 13856 21215 13890 21249
rect 13856 21147 13890 21181
rect 14852 23119 14886 23153
rect 14852 23051 14886 23085
rect 14852 22983 14886 23017
rect 14852 22915 14886 22949
rect 14852 22847 14886 22881
rect 14852 22779 14886 22813
rect 14852 22711 14886 22745
rect 14852 22643 14886 22677
rect 14852 22575 14886 22609
rect 14852 22507 14886 22541
rect 14852 22439 14886 22473
rect 14852 22371 14886 22405
rect 14852 22303 14886 22337
rect 14852 22235 14886 22269
rect 14852 22167 14886 22201
rect 14852 22099 14886 22133
rect 14852 22031 14886 22065
rect 14852 21963 14886 21997
rect 14852 21895 14886 21929
rect 14852 21827 14886 21861
rect 14852 21759 14886 21793
rect 14852 21691 14886 21725
rect 14852 21623 14886 21657
rect 14852 21555 14886 21589
rect 14852 21487 14886 21521
rect 14852 21419 14886 21453
rect 14852 21351 14886 21385
rect 14852 21283 14886 21317
rect 14852 21215 14886 21249
rect 13856 21079 13890 21113
rect 14852 21147 14886 21181
rect 14852 21079 14886 21113
rect 13980 20976 14014 21010
rect 14048 20976 14082 21010
rect 14116 20976 14150 21010
rect 14184 20976 14218 21010
rect 14252 20976 14286 21010
rect 14320 20976 14354 21010
rect 14388 20976 14422 21010
rect 14456 20976 14490 21010
rect 14524 20976 14558 21010
rect 14592 20976 14626 21010
rect 14660 20976 14694 21010
rect 14728 20976 14762 21010
rect 15176 23215 15210 23249
rect 15176 23147 15210 23181
rect 15176 23079 15210 23113
rect 15176 23011 15210 23045
rect 15176 22943 15210 22977
rect 15176 22875 15210 22909
rect 15176 22807 15210 22841
rect 15176 22739 15210 22773
rect 15176 22671 15210 22705
rect 15176 22603 15210 22637
rect 15176 22535 15210 22569
rect 15176 22467 15210 22501
rect 15176 22399 15210 22433
rect 15176 22331 15210 22365
rect 15176 22263 15210 22297
rect 15176 22195 15210 22229
rect 15176 22127 15210 22161
rect 15176 22059 15210 22093
rect 15176 21991 15210 22025
rect 15176 21923 15210 21957
rect 15176 21855 15210 21889
rect 15176 21787 15210 21821
rect 15176 21719 15210 21753
rect 15176 21651 15210 21685
rect 15176 21583 15210 21617
rect 15176 21515 15210 21549
rect 15176 21447 15210 21481
rect 15176 21379 15210 21413
rect 15176 21311 15210 21345
rect 15176 21243 15210 21277
rect 15176 21175 15210 21209
rect 15176 21107 15210 21141
rect 15472 23215 15506 23249
rect 15472 23147 15506 23181
rect 15472 23079 15506 23113
rect 15472 23011 15506 23045
rect 15472 22943 15506 22977
rect 15472 22875 15506 22909
rect 15472 22807 15506 22841
rect 15472 22739 15506 22773
rect 15472 22671 15506 22705
rect 15472 22603 15506 22637
rect 15472 22535 15506 22569
rect 15472 22467 15506 22501
rect 15472 22399 15506 22433
rect 15472 22331 15506 22365
rect 15472 22263 15506 22297
rect 15472 22195 15506 22229
rect 15472 22127 15506 22161
rect 15472 22059 15506 22093
rect 15472 21991 15506 22025
rect 15472 21923 15506 21957
rect 15472 21855 15506 21889
rect 15472 21787 15506 21821
rect 15472 21719 15506 21753
rect 15472 21651 15506 21685
rect 15472 21583 15506 21617
rect 15472 21515 15506 21549
rect 15472 21447 15506 21481
rect 15472 21379 15506 21413
rect 15472 21311 15506 21345
rect 15472 21243 15506 21277
rect 15472 21175 15506 21209
rect 15472 21107 15506 21141
rect 15290 20996 15324 21030
rect 15358 20996 15392 21030
rect 16548 23329 16582 23363
rect 16548 23261 16582 23295
rect 16548 23193 16582 23227
rect 16548 23125 16582 23159
rect 16548 23057 16582 23091
rect 16548 22989 16582 23023
rect 16548 22921 16582 22955
rect 16548 22853 16582 22887
rect 16548 22785 16582 22819
rect 16548 22717 16582 22751
rect 16548 22649 16582 22683
rect 16548 22581 16582 22615
rect 16548 22513 16582 22547
rect 16548 22445 16582 22479
rect 16548 22377 16582 22411
rect 16548 22309 16582 22343
rect 16548 22241 16582 22275
rect 16548 22173 16582 22207
rect 16548 22105 16582 22139
rect 16548 22037 16582 22071
rect 17736 24009 17770 24043
rect 17736 23941 17770 23975
rect 17736 23873 17770 23907
rect 17736 23805 17770 23839
rect 17736 23737 17770 23771
rect 17736 23669 17770 23703
rect 17736 23601 17770 23635
rect 17736 23533 17770 23567
rect 17736 23465 17770 23499
rect 17736 23397 17770 23431
rect 17736 23329 17770 23363
rect 17736 23261 17770 23295
rect 17736 23193 17770 23227
rect 17736 23125 17770 23159
rect 17736 23057 17770 23091
rect 17736 22989 17770 23023
rect 17736 22921 17770 22955
rect 17736 22853 17770 22887
rect 17736 22785 17770 22819
rect 17736 22717 17770 22751
rect 17736 22649 17770 22683
rect 17736 22581 17770 22615
rect 17736 22513 17770 22547
rect 17736 22445 17770 22479
rect 17736 22377 17770 22411
rect 17736 22309 17770 22343
rect 17736 22241 17770 22275
rect 17736 22173 17770 22207
rect 17736 22105 17770 22139
rect 16548 21969 16582 22003
rect 17736 22037 17770 22071
rect 17736 21969 17770 22003
rect 16666 21866 16700 21900
rect 16734 21866 16768 21900
rect 16802 21866 16836 21900
rect 16870 21866 16904 21900
rect 16938 21866 16972 21900
rect 17006 21866 17040 21900
rect 17074 21866 17108 21900
rect 17142 21866 17176 21900
rect 17210 21866 17244 21900
rect 17278 21866 17312 21900
rect 17346 21866 17380 21900
rect 17414 21866 17448 21900
rect 17482 21866 17516 21900
rect 17550 21866 17584 21900
rect 17618 21866 17652 21900
rect 16770 21446 16804 21480
rect 16838 21446 16872 21480
rect 16656 21325 16690 21359
rect 16656 21257 16690 21291
rect 16656 21189 16690 21223
rect 16656 21121 16690 21155
rect 16656 21053 16690 21087
rect 16656 20985 16690 21019
rect 16656 20917 16690 20951
rect 16656 20849 16690 20883
rect 16656 20781 16690 20815
rect 16656 20713 16690 20747
rect 16656 20645 16690 20679
rect 14826 20586 14860 20620
rect 14894 20586 14928 20620
rect 14962 20586 14996 20620
rect 15030 20586 15064 20620
rect 15098 20586 15132 20620
rect 15166 20586 15200 20620
rect 15234 20586 15268 20620
rect 15302 20586 15336 20620
rect 15370 20586 15404 20620
rect 15438 20586 15472 20620
rect 15506 20586 15540 20620
rect 14716 20466 14750 20500
rect 15616 20466 15650 20500
rect 14716 20398 14750 20432
rect 14716 20330 14750 20364
rect 14716 20262 14750 20296
rect 14716 20194 14750 20228
rect 14716 20126 14750 20160
rect 14716 20058 14750 20092
rect 14716 19990 14750 20024
rect 14716 19922 14750 19956
rect 13286 19826 13320 19860
rect 13354 19826 13388 19860
rect 13422 19826 13456 19860
rect 13490 19826 13524 19860
rect 13558 19826 13592 19860
rect 13626 19826 13660 19860
rect 13694 19826 13728 19860
rect 13762 19826 13796 19860
rect 13830 19826 13864 19860
rect 13898 19826 13932 19860
rect 13966 19826 14000 19860
rect 14034 19826 14068 19860
rect 14102 19826 14136 19860
rect 14170 19826 14204 19860
rect 14238 19826 14272 19860
rect 14306 19826 14340 19860
rect 13182 19721 13216 19755
rect 13182 19653 13216 19687
rect 13182 19585 13216 19619
rect 14410 19721 14444 19755
rect 14410 19653 14444 19687
rect 13182 19517 13216 19551
rect 13182 19449 13216 19483
rect 13182 19381 13216 19415
rect 13182 19313 13216 19347
rect 14410 19585 14444 19619
rect 14410 19517 14444 19551
rect 14410 19449 14444 19483
rect 14410 19381 14444 19415
rect 13182 19245 13216 19279
rect 13182 19177 13216 19211
rect 14410 19313 14444 19347
rect 14410 19245 14444 19279
rect 13182 19109 13216 19143
rect 13182 19041 13216 19075
rect 13182 18973 13216 19007
rect 14410 19177 14444 19211
rect 14410 19109 14444 19143
rect 14410 19041 14444 19075
rect 14410 18973 14444 19007
rect 14716 19854 14750 19888
rect 14716 19786 14750 19820
rect 14716 19718 14750 19752
rect 14716 19650 14750 19684
rect 14716 19582 14750 19616
rect 14716 19514 14750 19548
rect 14716 19446 14750 19480
rect 14716 19378 14750 19412
rect 14716 19310 14750 19344
rect 14716 19242 14750 19276
rect 14716 19174 14750 19208
rect 15616 20398 15650 20432
rect 15616 20330 15650 20364
rect 15616 20262 15650 20296
rect 15616 20194 15650 20228
rect 15616 20126 15650 20160
rect 16656 20577 16690 20611
rect 16656 20509 16690 20543
rect 16656 20441 16690 20475
rect 16656 20373 16690 20407
rect 16656 20305 16690 20339
rect 16656 20237 16690 20271
rect 16656 20169 16690 20203
rect 15616 20058 15650 20092
rect 15616 19990 15650 20024
rect 15616 19922 15650 19956
rect 15616 19854 15650 19888
rect 15616 19786 15650 19820
rect 15616 19718 15650 19752
rect 15616 19650 15650 19684
rect 15616 19582 15650 19616
rect 15616 19514 15650 19548
rect 15616 19446 15650 19480
rect 15616 19378 15650 19412
rect 15616 19310 15650 19344
rect 15616 19242 15650 19276
rect 15616 19174 15650 19208
rect 14716 19106 14750 19140
rect 15616 19106 15650 19140
rect 14826 18986 14860 19020
rect 14894 18986 14928 19020
rect 14962 18986 14996 19020
rect 15030 18986 15064 19020
rect 15098 18986 15132 19020
rect 15166 18986 15200 19020
rect 15234 18986 15268 19020
rect 15302 18986 15336 19020
rect 15370 18986 15404 19020
rect 15438 18986 15472 19020
rect 15506 18986 15540 19020
rect 15998 20100 16032 20134
rect 16066 20100 16100 20134
rect 16134 20100 16168 20134
rect 16202 20100 16236 20134
rect 16270 20100 16304 20134
rect 15876 19985 15910 20019
rect 16392 19985 16426 20019
rect 15876 19917 15910 19951
rect 15876 19849 15910 19883
rect 15876 19781 15910 19815
rect 15876 19713 15910 19747
rect 15876 19645 15910 19679
rect 15876 19577 15910 19611
rect 15876 19509 15910 19543
rect 15876 19441 15910 19475
rect 15876 19373 15910 19407
rect 15876 19305 15910 19339
rect 15876 19237 15910 19271
rect 15876 19169 15910 19203
rect 16392 19917 16426 19951
rect 16392 19849 16426 19883
rect 16392 19781 16426 19815
rect 16392 19713 16426 19747
rect 16392 19645 16426 19679
rect 16392 19577 16426 19611
rect 16392 19509 16426 19543
rect 16392 19441 16426 19475
rect 16392 19373 16426 19407
rect 16392 19305 16426 19339
rect 16392 19237 16426 19271
rect 16392 19169 16426 19203
rect 15876 19101 15910 19135
rect 16392 19101 16426 19135
rect 15998 18986 16032 19020
rect 16066 18986 16100 19020
rect 16134 18986 16168 19020
rect 16202 18986 16236 19020
rect 16270 18986 16304 19020
rect 16656 20101 16690 20135
rect 16656 20033 16690 20067
rect 16656 19965 16690 19999
rect 16656 19897 16690 19931
rect 16656 19829 16690 19863
rect 16656 19761 16690 19795
rect 16656 19693 16690 19727
rect 16656 19625 16690 19659
rect 16656 19557 16690 19591
rect 16656 19489 16690 19523
rect 16656 19421 16690 19455
rect 16656 19353 16690 19387
rect 16656 19285 16690 19319
rect 16656 19217 16690 19251
rect 16656 19149 16690 19183
rect 16656 19081 16690 19115
rect 16656 19013 16690 19047
rect 13182 18905 13216 18939
rect 13182 18837 13216 18871
rect 14410 18905 14444 18939
rect 14410 18837 14444 18871
rect 13182 18769 13216 18803
rect 13182 18701 13216 18735
rect 13182 18633 13216 18667
rect 13182 18565 13216 18599
rect 14410 18769 14444 18803
rect 16656 18945 16690 18979
rect 16656 18877 16690 18911
rect 16952 21325 16986 21359
rect 16952 21257 16986 21291
rect 16952 21189 16986 21223
rect 16952 21121 16986 21155
rect 16952 21053 16986 21087
rect 16952 20985 16986 21019
rect 16952 20917 16986 20951
rect 16952 20849 16986 20883
rect 16952 20781 16986 20815
rect 16952 20713 16986 20747
rect 16952 20645 16986 20679
rect 16952 20577 16986 20611
rect 16952 20509 16986 20543
rect 16952 20441 16986 20475
rect 16952 20373 16986 20407
rect 16952 20305 16986 20339
rect 16952 20237 16986 20271
rect 16952 20169 16986 20203
rect 16952 20101 16986 20135
rect 16952 20033 16986 20067
rect 16952 19965 16986 19999
rect 16952 19897 16986 19931
rect 16952 19829 16986 19863
rect 16952 19761 16986 19795
rect 16952 19693 16986 19727
rect 16952 19625 16986 19659
rect 16952 19557 16986 19591
rect 16952 19489 16986 19523
rect 16952 19421 16986 19455
rect 16952 19353 16986 19387
rect 16952 19285 16986 19319
rect 16952 19217 16986 19251
rect 16952 19149 16986 19183
rect 16952 19081 16986 19115
rect 16952 19013 16986 19047
rect 16952 18945 16986 18979
rect 16952 18877 16986 18911
rect 16770 18756 16804 18790
rect 16838 18756 16872 18790
rect 17380 21466 17414 21500
rect 17448 21466 17482 21500
rect 17266 21359 17300 21393
rect 17266 21291 17300 21325
rect 17266 21223 17300 21257
rect 17266 21155 17300 21189
rect 17266 21087 17300 21121
rect 17266 21019 17300 21053
rect 17266 20951 17300 20985
rect 17266 20883 17300 20917
rect 17266 20815 17300 20849
rect 17266 20747 17300 20781
rect 17266 20679 17300 20713
rect 17266 20611 17300 20645
rect 17266 20543 17300 20577
rect 17266 20475 17300 20509
rect 17266 20407 17300 20441
rect 17266 20339 17300 20373
rect 17266 20271 17300 20305
rect 17266 20203 17300 20237
rect 17266 20135 17300 20169
rect 17266 20067 17300 20101
rect 17266 19999 17300 20033
rect 17266 19931 17300 19965
rect 17266 19863 17300 19897
rect 17266 19795 17300 19829
rect 17266 19727 17300 19761
rect 17266 19659 17300 19693
rect 17266 19591 17300 19625
rect 17266 19523 17300 19557
rect 17266 19455 17300 19489
rect 17266 19387 17300 19421
rect 17266 19319 17300 19353
rect 17266 19251 17300 19285
rect 17266 19183 17300 19217
rect 17266 19115 17300 19149
rect 17266 19047 17300 19081
rect 17266 18979 17300 19013
rect 17266 18911 17300 18945
rect 17266 18843 17300 18877
rect 17266 18775 17300 18809
rect 14410 18701 14444 18735
rect 17266 18707 17300 18741
rect 14410 18633 14444 18667
rect 13182 18497 13216 18531
rect 13182 18429 13216 18463
rect 14410 18565 14444 18599
rect 14410 18497 14444 18531
rect 13182 18361 13216 18395
rect 13182 18293 13216 18327
rect 13182 18225 13216 18259
rect 13182 18157 13216 18191
rect 14410 18429 14444 18463
rect 14410 18361 14444 18395
rect 14410 18293 14444 18327
rect 14410 18225 14444 18259
rect 13182 18089 13216 18123
rect 13182 18021 13216 18055
rect 14410 18157 14444 18191
rect 14410 18089 14444 18123
rect 13182 17953 13216 17987
rect 13182 17885 13216 17919
rect 13182 17817 13216 17851
rect 14410 18021 14444 18055
rect 14410 17953 14444 17987
rect 15026 18634 15060 18668
rect 15094 18634 15128 18668
rect 14902 18513 14936 18547
rect 15218 18513 15252 18547
rect 14902 18445 14936 18479
rect 14902 18377 14936 18411
rect 14902 18309 14936 18343
rect 14902 18241 14936 18275
rect 14902 18173 14936 18207
rect 14902 18105 14936 18139
rect 14902 18037 14936 18071
rect 14410 17885 14444 17919
rect 14410 17817 14444 17851
rect 13182 17749 13216 17783
rect 13182 17681 13216 17715
rect 14410 17749 14444 17783
rect 14410 17681 14444 17715
rect 13182 17613 13216 17647
rect 13182 17545 13216 17579
rect 13182 17477 13216 17511
rect 13182 17409 13216 17443
rect 14410 17613 14444 17647
rect 14410 17545 14444 17579
rect 14410 17477 14444 17511
rect 13182 17341 13216 17375
rect 13182 17273 13216 17307
rect 14410 17409 14444 17443
rect 14410 17341 14444 17375
rect 13182 17205 13216 17239
rect 13182 17137 13216 17171
rect 13182 17069 13216 17103
rect 13182 17001 13216 17035
rect 14410 17273 14444 17307
rect 14410 17205 14444 17239
rect 14410 17137 14444 17171
rect 14410 17069 14444 17103
rect 13182 16933 13216 16967
rect 13182 16865 13216 16899
rect 14410 17001 14444 17035
rect 14410 16933 14444 16967
rect 14410 16865 14444 16899
rect 13286 16760 13320 16794
rect 13354 16760 13388 16794
rect 13422 16760 13456 16794
rect 13490 16760 13524 16794
rect 13558 16760 13592 16794
rect 13626 16760 13660 16794
rect 13694 16760 13728 16794
rect 13762 16760 13796 16794
rect 13830 16760 13864 16794
rect 13898 16760 13932 16794
rect 13966 16760 14000 16794
rect 14034 16760 14068 16794
rect 14102 16760 14136 16794
rect 14170 16760 14204 16794
rect 14238 16760 14272 16794
rect 14306 16760 14340 16794
rect 14626 17950 14660 17984
rect 14694 17950 14728 17984
rect 14512 17831 14546 17865
rect 14512 17763 14546 17797
rect 14512 17695 14546 17729
rect 14512 17627 14546 17661
rect 14512 17559 14546 17593
rect 14512 17491 14546 17525
rect 14512 17423 14546 17457
rect 14512 17355 14546 17389
rect 14512 17287 14546 17321
rect 14512 17219 14546 17253
rect 14512 17151 14546 17185
rect 14512 17083 14546 17117
rect 14512 17015 14546 17049
rect 14512 16947 14546 16981
rect 14512 16879 14546 16913
rect 14808 17831 14842 17865
rect 14808 17763 14842 17797
rect 14808 17695 14842 17729
rect 14808 17627 14842 17661
rect 14808 17559 14842 17593
rect 14808 17491 14842 17525
rect 14808 17423 14842 17457
rect 14808 17355 14842 17389
rect 14808 17287 14842 17321
rect 14808 17219 14842 17253
rect 14808 17151 14842 17185
rect 14808 17083 14842 17117
rect 14808 17015 14842 17049
rect 14808 16947 14842 16981
rect 14808 16879 14842 16913
rect 14626 16760 14660 16794
rect 14694 16760 14728 16794
rect 14902 17969 14936 18003
rect 14902 17901 14936 17935
rect 14902 17833 14936 17867
rect 14902 17765 14936 17799
rect 14902 17697 14936 17731
rect 14902 17629 14936 17663
rect 14902 17561 14936 17595
rect 14902 17493 14936 17527
rect 14902 17425 14936 17459
rect 14902 17357 14936 17391
rect 14902 17289 14936 17323
rect 14902 17221 14936 17255
rect 14902 17153 14936 17187
rect 14902 17085 14936 17119
rect 14902 17017 14936 17051
rect 14902 16949 14936 16983
rect 15218 18445 15252 18479
rect 15218 18377 15252 18411
rect 15218 18309 15252 18343
rect 15218 18241 15252 18275
rect 15218 18173 15252 18207
rect 15218 18105 15252 18139
rect 15218 18037 15252 18071
rect 15218 17969 15252 18003
rect 15218 17901 15252 17935
rect 15218 17833 15252 17867
rect 15218 17765 15252 17799
rect 15218 17697 15252 17731
rect 15218 17629 15252 17663
rect 15218 17561 15252 17595
rect 15218 17493 15252 17527
rect 15218 17425 15252 17459
rect 15218 17357 15252 17391
rect 15218 17289 15252 17323
rect 15218 17221 15252 17255
rect 15218 17153 15252 17187
rect 15218 17085 15252 17119
rect 15218 17017 15252 17051
rect 15218 16949 15252 16983
rect 14902 16881 14936 16915
rect 15218 16881 15252 16915
rect 15026 16760 15060 16794
rect 15094 16760 15128 16794
rect 15436 18634 15470 18668
rect 15504 18634 15538 18668
rect 15312 18513 15346 18547
rect 15628 18513 15662 18547
rect 15312 18445 15346 18479
rect 15312 18377 15346 18411
rect 15312 18309 15346 18343
rect 15312 18241 15346 18275
rect 15312 18173 15346 18207
rect 15312 18105 15346 18139
rect 15312 18037 15346 18071
rect 15312 17969 15346 18003
rect 15312 17901 15346 17935
rect 15312 17833 15346 17867
rect 15312 17765 15346 17799
rect 15312 17697 15346 17731
rect 15312 17629 15346 17663
rect 15312 17561 15346 17595
rect 15312 17493 15346 17527
rect 15312 17425 15346 17459
rect 15312 17357 15346 17391
rect 15312 17289 15346 17323
rect 15312 17221 15346 17255
rect 15312 17153 15346 17187
rect 15312 17085 15346 17119
rect 15312 17017 15346 17051
rect 15312 16949 15346 16983
rect 15628 18445 15662 18479
rect 15628 18377 15662 18411
rect 15628 18309 15662 18343
rect 15628 18241 15662 18275
rect 15628 18173 15662 18207
rect 15628 18105 15662 18139
rect 15628 18037 15662 18071
rect 15628 17969 15662 18003
rect 16238 18651 16272 18685
rect 16306 18651 16340 18685
rect 16124 18522 16158 18556
rect 16124 18454 16158 18488
rect 16124 18386 16158 18420
rect 16124 18318 16158 18352
rect 16124 18250 16158 18284
rect 16124 18182 16158 18216
rect 16124 18114 16158 18148
rect 16124 18046 16158 18080
rect 15628 17901 15662 17935
rect 15628 17833 15662 17867
rect 15628 17765 15662 17799
rect 15628 17697 15662 17731
rect 15628 17629 15662 17663
rect 15628 17561 15662 17595
rect 15628 17493 15662 17527
rect 15628 17425 15662 17459
rect 15628 17357 15662 17391
rect 15628 17289 15662 17323
rect 15628 17221 15662 17255
rect 15628 17153 15662 17187
rect 15628 17085 15662 17119
rect 15628 17017 15662 17051
rect 15628 16949 15662 16983
rect 15312 16881 15346 16915
rect 15628 16881 15662 16915
rect 15436 16760 15470 16794
rect 15504 16760 15538 16794
rect 15846 17950 15880 17984
rect 15914 17950 15948 17984
rect 15732 17831 15766 17865
rect 15732 17763 15766 17797
rect 15732 17695 15766 17729
rect 15732 17627 15766 17661
rect 15732 17559 15766 17593
rect 15732 17491 15766 17525
rect 15732 17423 15766 17457
rect 15732 17355 15766 17389
rect 15732 17287 15766 17321
rect 15732 17219 15766 17253
rect 15732 17151 15766 17185
rect 15732 17083 15766 17117
rect 15732 17015 15766 17049
rect 15732 16947 15766 16981
rect 15732 16879 15766 16913
rect 16028 17831 16062 17865
rect 16028 17763 16062 17797
rect 16028 17695 16062 17729
rect 16028 17627 16062 17661
rect 16028 17559 16062 17593
rect 16028 17491 16062 17525
rect 16028 17423 16062 17457
rect 16028 17355 16062 17389
rect 16028 17287 16062 17321
rect 16028 17219 16062 17253
rect 16028 17151 16062 17185
rect 16028 17083 16062 17117
rect 16028 17015 16062 17049
rect 16028 16947 16062 16981
rect 16028 16879 16062 16913
rect 15846 16760 15880 16794
rect 15914 16760 15948 16794
rect 16124 17978 16158 18012
rect 16124 17910 16158 17944
rect 16124 17842 16158 17876
rect 16124 17774 16158 17808
rect 16124 17706 16158 17740
rect 16124 17638 16158 17672
rect 16124 17570 16158 17604
rect 16124 17502 16158 17536
rect 16124 17434 16158 17468
rect 16124 17366 16158 17400
rect 16124 17298 16158 17332
rect 16124 17230 16158 17264
rect 16124 17162 16158 17196
rect 16124 17094 16158 17128
rect 16124 17026 16158 17060
rect 16124 16958 16158 16992
rect 16124 16890 16158 16924
rect 16420 18522 16454 18556
rect 16420 18454 16454 18488
rect 17266 18639 17300 18673
rect 17266 18571 17300 18605
rect 17266 18503 17300 18537
rect 16420 18386 16454 18420
rect 16420 18318 16454 18352
rect 16420 18250 16454 18284
rect 16420 18182 16454 18216
rect 16782 18426 16816 18460
rect 16850 18426 16884 18460
rect 16686 18330 16720 18364
rect 16686 18262 16720 18296
rect 16946 18330 16980 18364
rect 16946 18262 16980 18296
rect 16782 18166 16816 18200
rect 16850 18166 16884 18200
rect 17266 18435 17300 18469
rect 17266 18367 17300 18401
rect 17266 18299 17300 18333
rect 17266 18231 17300 18265
rect 16420 18114 16454 18148
rect 16420 18046 16454 18080
rect 16420 17978 16454 18012
rect 16420 17910 16454 17944
rect 16420 17842 16454 17876
rect 16420 17774 16454 17808
rect 16420 17706 16454 17740
rect 16420 17638 16454 17672
rect 16420 17570 16454 17604
rect 16420 17502 16454 17536
rect 16420 17434 16454 17468
rect 16420 17366 16454 17400
rect 17266 18163 17300 18197
rect 17266 18095 17300 18129
rect 17266 18027 17300 18061
rect 17266 17959 17300 17993
rect 17266 17891 17300 17925
rect 17266 17823 17300 17857
rect 17266 17755 17300 17789
rect 17266 17687 17300 17721
rect 17266 17619 17300 17653
rect 17266 17551 17300 17585
rect 17266 17483 17300 17517
rect 17562 21359 17596 21393
rect 17562 21291 17596 21325
rect 17562 21223 17596 21257
rect 17562 21155 17596 21189
rect 17562 21087 17596 21121
rect 17562 21019 17596 21053
rect 17562 20951 17596 20985
rect 17562 20883 17596 20917
rect 17562 20815 17596 20849
rect 17562 20747 17596 20781
rect 17562 20679 17596 20713
rect 17562 20611 17596 20645
rect 17562 20543 17596 20577
rect 17562 20475 17596 20509
rect 17562 20407 17596 20441
rect 17562 20339 17596 20373
rect 17562 20271 17596 20305
rect 17562 20203 17596 20237
rect 17562 20135 17596 20169
rect 17562 20067 17596 20101
rect 17562 19999 17596 20033
rect 17562 19931 17596 19965
rect 17562 19863 17596 19897
rect 17562 19795 17596 19829
rect 17562 19727 17596 19761
rect 17562 19659 17596 19693
rect 17562 19591 17596 19625
rect 17562 19523 17596 19557
rect 17562 19455 17596 19489
rect 17562 19387 17596 19421
rect 17562 19319 17596 19353
rect 17562 19251 17596 19285
rect 17562 19183 17596 19217
rect 17562 19115 17596 19149
rect 17562 19047 17596 19081
rect 17562 18979 17596 19013
rect 17562 18911 17596 18945
rect 17562 18843 17596 18877
rect 17562 18775 17596 18809
rect 17562 18707 17596 18741
rect 17562 18639 17596 18673
rect 17562 18571 17596 18605
rect 17562 18503 17596 18537
rect 17562 18435 17596 18469
rect 17562 18367 17596 18401
rect 17562 18299 17596 18333
rect 17562 18231 17596 18265
rect 17562 18163 17596 18197
rect 17562 18095 17596 18129
rect 17562 18027 17596 18061
rect 17562 17959 17596 17993
rect 17562 17891 17596 17925
rect 17562 17823 17596 17857
rect 17562 17755 17596 17789
rect 17562 17687 17596 17721
rect 17562 17619 17596 17653
rect 17562 17551 17596 17585
rect 17562 17483 17596 17517
rect 17380 17376 17414 17410
rect 17448 17376 17482 17410
rect 16420 17298 16454 17332
rect 16420 17230 16454 17264
rect 16420 17162 16454 17196
rect 16420 17094 16454 17128
rect 16420 17026 16454 17060
rect 16420 16958 16454 16992
rect 16420 16890 16454 16924
rect 16238 16761 16272 16795
rect 16306 16761 16340 16795
rect 14432 16044 14466 16078
rect 14500 16044 14534 16078
rect 14568 16044 14602 16078
rect 14636 16044 14670 16078
rect 14704 16044 14738 16078
rect 14772 16044 14806 16078
rect 14840 16044 14874 16078
rect 14908 16044 14942 16078
rect 14976 16044 15010 16078
rect 15044 16044 15078 16078
rect 15112 16044 15146 16078
rect 15180 16044 15214 16078
rect 14308 15941 14342 15975
rect 14308 15873 14342 15907
rect 15304 15941 15338 15975
rect 14308 15805 14342 15839
rect 14308 15737 14342 15771
rect 14308 15669 14342 15703
rect 13582 15604 13616 15638
rect 13650 15604 13684 15638
rect 13458 15483 13492 15517
rect 13774 15483 13808 15517
rect 13458 15415 13492 15449
rect 13458 15347 13492 15381
rect 13458 15279 13492 15313
rect 13458 15211 13492 15245
rect 13458 15143 13492 15177
rect 13458 15075 13492 15109
rect 13458 15007 13492 15041
rect 13458 14939 13492 14973
rect 13458 14871 13492 14905
rect 13458 14803 13492 14837
rect 13458 14735 13492 14769
rect 13458 14667 13492 14701
rect 13458 14599 13492 14633
rect 13458 14531 13492 14565
rect 13458 14463 13492 14497
rect 13458 14395 13492 14429
rect 13458 14327 13492 14361
rect 13458 14259 13492 14293
rect 13458 14191 13492 14225
rect 13458 14123 13492 14157
rect 13458 14055 13492 14089
rect 13458 13987 13492 14021
rect 13458 13919 13492 13953
rect 13774 15415 13808 15449
rect 13774 15347 13808 15381
rect 13774 15279 13808 15313
rect 13774 15211 13808 15245
rect 13774 15143 13808 15177
rect 13774 15075 13808 15109
rect 13774 15007 13808 15041
rect 13774 14939 13808 14973
rect 13774 14871 13808 14905
rect 13774 14803 13808 14837
rect 13774 14735 13808 14769
rect 13774 14667 13808 14701
rect 13774 14599 13808 14633
rect 13774 14531 13808 14565
rect 13774 14463 13808 14497
rect 13774 14395 13808 14429
rect 13774 14327 13808 14361
rect 13774 14259 13808 14293
rect 13774 14191 13808 14225
rect 13774 14123 13808 14157
rect 13774 14055 13808 14089
rect 13774 13987 13808 14021
rect 13774 13919 13808 13953
rect 13458 13851 13492 13885
rect 13774 13851 13808 13885
rect 13582 13730 13616 13764
rect 13650 13730 13684 13764
rect 14308 15601 14342 15635
rect 14308 15533 14342 15567
rect 14308 15465 14342 15499
rect 14308 15397 14342 15431
rect 14308 15329 14342 15363
rect 14308 15261 14342 15295
rect 14308 15193 14342 15227
rect 14308 15125 14342 15159
rect 14308 15057 14342 15091
rect 14308 14989 14342 15023
rect 14308 14921 14342 14955
rect 14308 14853 14342 14887
rect 14308 14785 14342 14819
rect 14308 14717 14342 14751
rect 14308 14649 14342 14683
rect 14308 14581 14342 14615
rect 14308 14513 14342 14547
rect 14308 14445 14342 14479
rect 14308 14377 14342 14411
rect 14308 14309 14342 14343
rect 14308 14241 14342 14275
rect 14308 14173 14342 14207
rect 14308 14105 14342 14139
rect 14308 14037 14342 14071
rect 14308 13969 14342 14003
rect 14308 13901 14342 13935
rect 15304 15873 15338 15907
rect 15304 15805 15338 15839
rect 15304 15737 15338 15771
rect 15304 15669 15338 15703
rect 15304 15601 15338 15635
rect 15304 15533 15338 15567
rect 15304 15465 15338 15499
rect 15304 15397 15338 15431
rect 15304 15329 15338 15363
rect 15304 15261 15338 15295
rect 15304 15193 15338 15227
rect 15304 15125 15338 15159
rect 15304 15057 15338 15091
rect 15304 14989 15338 15023
rect 15304 14921 15338 14955
rect 15304 14853 15338 14887
rect 15304 14785 15338 14819
rect 15304 14717 15338 14751
rect 15304 14649 15338 14683
rect 15304 14581 15338 14615
rect 15304 14513 15338 14547
rect 15304 14445 15338 14479
rect 15304 14377 15338 14411
rect 15304 14309 15338 14343
rect 15304 14241 15338 14275
rect 15304 14173 15338 14207
rect 15304 14105 15338 14139
rect 15304 14037 15338 14071
rect 15304 13969 15338 14003
rect 14308 13833 14342 13867
rect 15304 13901 15338 13935
rect 15304 13833 15338 13867
rect 14432 13730 14466 13764
rect 14500 13730 14534 13764
rect 14568 13730 14602 13764
rect 14636 13730 14670 13764
rect 14704 13730 14738 13764
rect 14772 13730 14806 13764
rect 14840 13730 14874 13764
rect 14908 13730 14942 13764
rect 14976 13730 15010 13764
rect 15044 13730 15078 13764
rect 15112 13730 15146 13764
rect 15180 13730 15214 13764
rect 16132 16060 16166 16094
rect 16200 16060 16234 16094
rect 16018 15949 16052 15983
rect 16018 15881 16052 15915
rect 16018 15813 16052 15847
rect 16018 15745 16052 15779
rect 16018 15677 16052 15711
rect 16018 15609 16052 15643
rect 16018 15541 16052 15575
rect 16018 15473 16052 15507
rect 16018 15405 16052 15439
rect 16018 15337 16052 15371
rect 16018 15269 16052 15303
rect 16018 15201 16052 15235
rect 16018 15133 16052 15167
rect 16018 15065 16052 15099
rect 16018 14997 16052 15031
rect 16018 14929 16052 14963
rect 16018 14861 16052 14895
rect 16018 14793 16052 14827
rect 16018 14725 16052 14759
rect 16018 14657 16052 14691
rect 16018 14589 16052 14623
rect 16018 14521 16052 14555
rect 16018 14453 16052 14487
rect 16018 14385 16052 14419
rect 16018 14317 16052 14351
rect 16018 14249 16052 14283
rect 16018 14181 16052 14215
rect 16018 14113 16052 14147
rect 16018 14045 16052 14079
rect 16018 13977 16052 14011
rect 16018 13909 16052 13943
rect 16018 13841 16052 13875
rect 16314 15949 16348 15983
rect 16314 15881 16348 15915
rect 16314 15813 16348 15847
rect 16314 15745 16348 15779
rect 16314 15677 16348 15711
rect 16314 15609 16348 15643
rect 16314 15541 16348 15575
rect 16314 15473 16348 15507
rect 16314 15405 16348 15439
rect 16314 15337 16348 15371
rect 16314 15269 16348 15303
rect 16314 15201 16348 15235
rect 16314 15133 16348 15167
rect 16314 15065 16348 15099
rect 16314 14997 16348 15031
rect 16314 14929 16348 14963
rect 16314 14861 16348 14895
rect 16314 14793 16348 14827
rect 16314 14725 16348 14759
rect 16314 14657 16348 14691
rect 16314 14589 16348 14623
rect 16314 14521 16348 14555
rect 16314 14453 16348 14487
rect 16314 14385 16348 14419
rect 16314 14317 16348 14351
rect 16314 14249 16348 14283
rect 16314 14181 16348 14215
rect 16314 14113 16348 14147
rect 16314 14045 16348 14079
rect 16314 13977 16348 14011
rect 16314 13909 16348 13943
rect 16314 13841 16348 13875
rect 16132 13730 16166 13764
rect 16200 13730 16234 13764
rect 13329 13512 13363 13546
rect 13397 13512 13431 13546
rect 13465 13512 13499 13546
rect 13533 13512 13567 13546
rect 13601 13512 13635 13546
rect 13669 13512 13703 13546
rect 13737 13512 13771 13546
rect 13805 13512 13839 13546
rect 13873 13512 13907 13546
rect 13941 13512 13975 13546
rect 14009 13512 14043 13546
rect 14077 13512 14111 13546
rect 14145 13512 14179 13546
rect 14213 13512 14247 13546
rect 14281 13512 14315 13546
rect 14349 13512 14383 13546
rect 14417 13512 14451 13546
rect 14485 13512 14519 13546
rect 14553 13512 14587 13546
rect 14621 13512 14655 13546
rect 14689 13512 14723 13546
rect 14757 13512 14791 13546
rect 14825 13512 14859 13546
rect 14893 13512 14927 13546
rect 14961 13512 14995 13546
rect 15029 13512 15063 13546
rect 15097 13512 15131 13546
rect 15165 13512 15199 13546
rect 15233 13512 15267 13546
rect 15301 13512 15335 13546
rect 15369 13512 15403 13546
rect 15437 13512 15471 13546
rect 15505 13512 15539 13546
rect 15573 13512 15607 13546
rect 15641 13512 15675 13546
rect 15709 13512 15743 13546
rect 15777 13512 15811 13546
rect 15845 13512 15879 13546
rect 15913 13512 15947 13546
rect 15981 13512 16015 13546
rect 16049 13512 16083 13546
rect 16117 13512 16151 13546
rect 16185 13512 16219 13546
rect 16253 13512 16287 13546
rect 16321 13512 16355 13546
rect 16389 13512 16423 13546
rect 16457 13512 16491 13546
rect 16525 13512 16559 13546
rect 16593 13512 16627 13546
rect 16661 13512 16695 13546
rect 16729 13512 16763 13546
rect 16797 13512 16831 13546
rect 16865 13512 16899 13546
rect 16933 13512 16967 13546
rect 17001 13512 17035 13546
rect 17069 13512 17103 13546
rect 17137 13512 17171 13546
rect 17205 13512 17239 13546
rect 17273 13512 17307 13546
rect 17341 13512 17375 13546
rect 17409 13512 17443 13546
rect 17477 13512 17511 13546
rect 17545 13512 17579 13546
rect 13122 13382 13156 13416
rect 13122 13314 13156 13348
rect 17785 13391 17819 13425
rect 13122 13246 13156 13280
rect 13122 13178 13156 13212
rect 13122 13110 13156 13144
rect 13122 13042 13156 13076
rect 17785 13323 17819 13357
rect 17785 13255 17819 13289
rect 17785 13187 17819 13221
rect 17785 13119 17819 13153
rect 13122 12974 13156 13008
rect 13122 12906 13156 12940
rect 13122 12838 13156 12872
rect 13122 12770 13156 12804
rect 13122 12702 13156 12736
rect 13122 12634 13156 12668
rect 13122 12566 13156 12600
rect 13122 12498 13156 12532
rect 13122 12430 13156 12464
rect 13122 12362 13156 12396
rect 13122 12294 13156 12328
rect 13122 12226 13156 12260
rect 13122 12158 13156 12192
rect 13122 12090 13156 12124
rect 13122 12022 13156 12056
rect 13122 11954 13156 11988
rect 13122 11886 13156 11920
rect 13122 11818 13156 11852
rect 13122 11750 13156 11784
rect 13122 11682 13156 11716
rect 13122 11614 13156 11648
rect 13122 11546 13156 11580
rect 13122 11478 13156 11512
rect 13122 11410 13156 11444
rect 13122 11342 13156 11376
rect 13122 11274 13156 11308
rect 13122 11206 13156 11240
rect 13122 11138 13156 11172
rect 13122 11070 13156 11104
rect 17785 13051 17819 13085
rect 17785 12983 17819 13017
rect 17785 12915 17819 12949
rect 17785 12847 17819 12881
rect 17785 12779 17819 12813
rect 17785 12711 17819 12745
rect 17785 12643 17819 12677
rect 17785 12575 17819 12609
rect 17785 12507 17819 12541
rect 17785 12439 17819 12473
rect 17785 12371 17819 12405
rect 17785 12303 17819 12337
rect 17785 12235 17819 12269
rect 17785 12167 17819 12201
rect 17785 12099 17819 12133
rect 17785 12031 17819 12065
rect 17785 11963 17819 11997
rect 17785 11895 17819 11929
rect 17785 11827 17819 11861
rect 17785 11759 17819 11793
rect 17785 11691 17819 11725
rect 17785 11623 17819 11657
rect 17785 11555 17819 11589
rect 17785 11487 17819 11521
rect 17785 11419 17819 11453
rect 17785 11351 17819 11385
rect 17785 11283 17819 11317
rect 17785 11215 17819 11249
rect 17785 11147 17819 11181
rect 17785 11079 17819 11113
rect 13122 11002 13156 11036
rect 13122 10934 13156 10968
rect 13122 10866 13156 10900
rect 17785 11011 17819 11045
rect 17785 10943 17819 10977
rect 13122 10798 13156 10832
rect 17785 10875 17819 10909
rect 17785 10807 17819 10841
rect 13371 10659 13405 10693
rect 13439 10659 13473 10693
rect 13507 10659 13541 10693
rect 13575 10659 13609 10693
rect 13643 10659 13677 10693
rect 13711 10659 13745 10693
rect 13779 10659 13813 10693
rect 13847 10659 13881 10693
rect 13915 10659 13949 10693
rect 13983 10659 14017 10693
rect 14051 10659 14085 10693
rect 14119 10659 14153 10693
rect 14187 10659 14221 10693
rect 14255 10659 14289 10693
rect 14323 10659 14357 10693
rect 14391 10659 14425 10693
rect 14459 10659 14493 10693
rect 14527 10659 14561 10693
rect 14595 10659 14629 10693
rect 14663 10659 14697 10693
rect 14731 10659 14765 10693
rect 14799 10659 14833 10693
rect 14867 10659 14901 10693
rect 14935 10659 14969 10693
rect 15003 10659 15037 10693
rect 15071 10659 15105 10693
rect 15139 10659 15173 10693
rect 15207 10659 15241 10693
rect 15275 10659 15309 10693
rect 15343 10659 15377 10693
rect 15411 10659 15445 10693
rect 15479 10659 15513 10693
rect 15547 10659 15581 10693
rect 15615 10659 15649 10693
rect 15683 10659 15717 10693
rect 15751 10659 15785 10693
rect 15819 10659 15853 10693
rect 15887 10659 15921 10693
rect 15955 10659 15989 10693
rect 16023 10659 16057 10693
rect 16091 10659 16125 10693
rect 16159 10659 16193 10693
rect 16227 10659 16261 10693
rect 16295 10659 16329 10693
rect 16363 10659 16397 10693
rect 16431 10659 16465 10693
rect 16499 10659 16533 10693
rect 16567 10659 16601 10693
rect 16635 10659 16669 10693
rect 16703 10659 16737 10693
rect 16771 10659 16805 10693
rect 16839 10659 16873 10693
rect 16907 10659 16941 10693
rect 16975 10659 17009 10693
rect 17043 10659 17077 10693
rect 17111 10659 17145 10693
rect 17179 10659 17213 10693
rect 17247 10659 17281 10693
rect 17315 10659 17349 10693
rect 17383 10659 17417 10693
rect 17451 10659 17485 10693
rect 17519 10659 17553 10693
rect 17587 10659 17621 10693
<< nsubdiffcont >>
rect 15838 23338 15872 23372
rect 15906 23338 15940 23372
rect 15974 23338 16008 23372
rect 16042 23338 16076 23372
rect 16110 23338 16144 23372
rect 15716 23226 15750 23260
rect 16232 23226 16266 23260
rect 15716 23158 15750 23192
rect 15716 23090 15750 23124
rect 15716 23022 15750 23056
rect 15716 22954 15750 22988
rect 15716 22886 15750 22920
rect 15716 22818 15750 22852
rect 15716 22750 15750 22784
rect 15716 22682 15750 22716
rect 15716 22614 15750 22648
rect 15716 22546 15750 22580
rect 15716 22478 15750 22512
rect 15716 22410 15750 22444
rect 15716 22342 15750 22376
rect 15716 22274 15750 22308
rect 15716 22206 15750 22240
rect 15716 22138 15750 22172
rect 15716 22070 15750 22104
rect 15716 22002 15750 22036
rect 15716 21934 15750 21968
rect 15716 21866 15750 21900
rect 15716 21798 15750 21832
rect 15716 21730 15750 21764
rect 15716 21662 15750 21696
rect 15716 21594 15750 21628
rect 15716 21526 15750 21560
rect 15716 21458 15750 21492
rect 15716 21390 15750 21424
rect 15716 21322 15750 21356
rect 15716 21254 15750 21288
rect 15716 21186 15750 21220
rect 16232 23158 16266 23192
rect 16232 23090 16266 23124
rect 16232 23022 16266 23056
rect 16232 22954 16266 22988
rect 16232 22886 16266 22920
rect 16232 22818 16266 22852
rect 16232 22750 16266 22784
rect 16232 22682 16266 22716
rect 16232 22614 16266 22648
rect 16232 22546 16266 22580
rect 16232 22478 16266 22512
rect 16232 22410 16266 22444
rect 16232 22342 16266 22376
rect 16232 22274 16266 22308
rect 16232 22206 16266 22240
rect 16232 22138 16266 22172
rect 16232 22070 16266 22104
rect 16232 22002 16266 22036
rect 16232 21934 16266 21968
rect 16232 21866 16266 21900
rect 16232 21798 16266 21832
rect 16232 21730 16266 21764
rect 16232 21662 16266 21696
rect 16232 21594 16266 21628
rect 16232 21526 16266 21560
rect 16232 21458 16266 21492
rect 16232 21390 16266 21424
rect 16232 21322 16266 21356
rect 16232 21254 16266 21288
rect 16232 21186 16266 21220
rect 15716 21118 15750 21152
rect 16232 21118 16266 21152
rect 15838 21006 15872 21040
rect 15906 21006 15940 21040
rect 15974 21006 16008 21040
rect 16042 21006 16076 21040
rect 16110 21006 16144 21040
rect 17100 16092 17134 16126
rect 17168 16092 17202 16126
rect 17236 16092 17270 16126
rect 17304 16092 17338 16126
rect 17372 16092 17406 16126
rect 16978 15980 17012 16014
rect 16978 15912 17012 15946
rect 17494 15980 17528 16014
rect 16978 15844 17012 15878
rect 16978 15776 17012 15810
rect 16978 15708 17012 15742
rect 16978 15640 17012 15674
rect 16978 15572 17012 15606
rect 16978 15504 17012 15538
rect 16978 15436 17012 15470
rect 16978 15368 17012 15402
rect 16978 15300 17012 15334
rect 16978 15232 17012 15266
rect 16978 15164 17012 15198
rect 16978 15096 17012 15130
rect 16978 15028 17012 15062
rect 16978 14960 17012 14994
rect 16978 14892 17012 14926
rect 16978 14824 17012 14858
rect 16978 14756 17012 14790
rect 16978 14688 17012 14722
rect 16978 14620 17012 14654
rect 16978 14552 17012 14586
rect 16978 14484 17012 14518
rect 16978 14416 17012 14450
rect 16978 14348 17012 14382
rect 16978 14280 17012 14314
rect 16978 14212 17012 14246
rect 16978 14144 17012 14178
rect 16978 14076 17012 14110
rect 16978 14008 17012 14042
rect 16978 13940 17012 13974
rect 17494 15912 17528 15946
rect 17494 15844 17528 15878
rect 17494 15776 17528 15810
rect 17494 15708 17528 15742
rect 17494 15640 17528 15674
rect 17494 15572 17528 15606
rect 17494 15504 17528 15538
rect 17494 15436 17528 15470
rect 17494 15368 17528 15402
rect 17494 15300 17528 15334
rect 17494 15232 17528 15266
rect 17494 15164 17528 15198
rect 17494 15096 17528 15130
rect 17494 15028 17528 15062
rect 17494 14960 17528 14994
rect 17494 14892 17528 14926
rect 17494 14824 17528 14858
rect 17494 14756 17528 14790
rect 17494 14688 17528 14722
rect 17494 14620 17528 14654
rect 17494 14552 17528 14586
rect 17494 14484 17528 14518
rect 17494 14416 17528 14450
rect 17494 14348 17528 14382
rect 17494 14280 17528 14314
rect 17494 14212 17528 14246
rect 17494 14144 17528 14178
rect 17494 14076 17528 14110
rect 17494 14008 17528 14042
rect 17494 13940 17528 13974
rect 16978 13872 17012 13906
rect 17494 13872 17528 13906
rect 17100 13760 17134 13794
rect 17168 13760 17202 13794
rect 17236 13760 17270 13794
rect 17304 13760 17338 13794
rect 17372 13760 17406 13794
<< poly >>
rect 16710 24112 16860 24130
rect 16710 24078 16806 24112
rect 16840 24078 16860 24112
rect 16710 24060 16860 24078
rect 16982 24112 17048 24128
rect 16982 24078 16998 24112
rect 17032 24078 17048 24112
rect 16712 24040 16742 24060
rect 16808 24040 16838 24060
rect 16904 24040 16934 24066
rect 16982 24062 17048 24078
rect 17174 24112 17240 24128
rect 17174 24078 17190 24112
rect 17224 24078 17240 24112
rect 17000 24040 17030 24062
rect 17096 24040 17126 24066
rect 17174 24062 17240 24078
rect 17366 24112 17432 24128
rect 17366 24078 17382 24112
rect 17416 24078 17432 24112
rect 17192 24040 17222 24062
rect 17288 24040 17318 24066
rect 17366 24062 17432 24078
rect 17558 24112 17624 24128
rect 17558 24078 17574 24112
rect 17608 24078 17624 24112
rect 17384 24040 17414 24062
rect 17480 24040 17510 24066
rect 17558 24062 17624 24078
rect 17576 24040 17606 24062
rect 14020 23222 14164 23238
rect 14020 23188 14114 23222
rect 14148 23188 14164 23222
rect 14020 23172 14164 23188
rect 14290 23222 14356 23238
rect 14290 23188 14306 23222
rect 14340 23188 14356 23222
rect 14020 23150 14050 23172
rect 14116 23150 14146 23172
rect 14212 23150 14242 23176
rect 14290 23172 14356 23188
rect 14482 23222 14548 23238
rect 14482 23188 14498 23222
rect 14532 23188 14548 23222
rect 14308 23150 14338 23172
rect 14404 23150 14434 23176
rect 14482 23172 14548 23188
rect 14674 23222 14740 23238
rect 14674 23188 14690 23222
rect 14724 23188 14740 23222
rect 14500 23150 14530 23172
rect 14596 23150 14626 23176
rect 14674 23172 14740 23188
rect 14692 23150 14722 23172
rect 14020 21128 14050 21150
rect 14002 21112 14068 21128
rect 14116 21124 14146 21150
rect 14212 21128 14242 21150
rect 14002 21078 14018 21112
rect 14052 21078 14068 21112
rect 14002 21062 14068 21078
rect 14194 21112 14260 21128
rect 14308 21124 14338 21150
rect 14404 21128 14434 21150
rect 14194 21078 14210 21112
rect 14244 21078 14260 21112
rect 14194 21062 14260 21078
rect 14386 21112 14452 21128
rect 14500 21124 14530 21150
rect 14596 21128 14626 21150
rect 14692 21128 14722 21150
rect 14386 21078 14402 21112
rect 14436 21078 14452 21112
rect 14386 21062 14452 21078
rect 14578 21112 14722 21128
rect 14578 21078 14594 21112
rect 14628 21078 14722 21112
rect 14578 21062 14722 21078
rect 15958 23270 16024 23286
rect 15958 23236 15974 23270
rect 16008 23236 16024 23270
rect 15958 23220 16024 23236
rect 15880 23189 15910 23215
rect 15976 23189 16006 23220
rect 16072 23189 16102 23215
rect 16712 22018 16742 22040
rect 16694 22002 16760 22018
rect 16808 22014 16838 22040
rect 16904 22018 16934 22040
rect 16694 21968 16710 22002
rect 16744 21968 16760 22002
rect 16694 21952 16760 21968
rect 16886 22002 16952 22018
rect 17000 22014 17030 22040
rect 17096 22018 17126 22040
rect 16886 21968 16902 22002
rect 16936 21968 16952 22002
rect 16886 21952 16952 21968
rect 17078 22002 17144 22018
rect 17192 22014 17222 22040
rect 17288 22018 17318 22040
rect 17078 21968 17094 22002
rect 17128 21968 17144 22002
rect 17078 21952 17144 21968
rect 17270 22002 17336 22018
rect 17384 22014 17414 22040
rect 17480 22020 17510 22040
rect 17576 22020 17606 22040
rect 17270 21968 17286 22002
rect 17320 21968 17336 22002
rect 17270 21952 17336 21968
rect 17460 22002 17610 22020
rect 17460 21968 17478 22002
rect 17512 21968 17610 22002
rect 17460 21950 17610 21968
rect 15880 21160 15910 21189
rect 15976 21160 16006 21189
rect 16072 21160 16102 21189
rect 15861 21142 16120 21160
rect 15861 21108 15878 21142
rect 15912 21108 16070 21142
rect 16104 21108 16120 21142
rect 15861 21091 16120 21108
rect 14880 20518 15490 20540
rect 14880 20484 14974 20518
rect 15008 20484 15166 20518
rect 15200 20484 15358 20518
rect 15392 20484 15490 20518
rect 14880 20470 15490 20484
rect 14880 20446 14910 20470
rect 14958 20468 15024 20470
rect 14976 20446 15006 20468
rect 15072 20446 15102 20470
rect 15150 20468 15216 20470
rect 15168 20446 15198 20468
rect 15264 20446 15294 20470
rect 15342 20468 15408 20470
rect 15360 20446 15390 20468
rect 15456 20446 15486 20470
rect 14880 19140 14910 19160
rect 14976 19140 15006 19160
rect 15072 19140 15102 19160
rect 15168 19140 15198 19160
rect 15264 19140 15294 19160
rect 15360 19140 15390 19160
rect 15456 19140 15486 19160
rect 14860 19122 15510 19140
rect 14860 19088 14878 19122
rect 14912 19088 15070 19122
rect 15104 19088 15262 19122
rect 15296 19088 15454 19122
rect 15488 19088 15510 19122
rect 14860 19070 15510 19088
rect 16040 20032 16270 20050
rect 16040 19998 16134 20032
rect 16168 19998 16270 20032
rect 16040 19980 16270 19998
rect 16040 19960 16070 19980
rect 16136 19960 16166 19980
rect 16232 19960 16262 19980
rect 16040 19140 16070 19160
rect 16136 19140 16166 19160
rect 16232 19140 16262 19160
rect 16020 19122 16280 19140
rect 16020 19088 16038 19122
rect 16072 19088 16230 19122
rect 16264 19088 16280 19122
rect 16020 19070 16280 19088
rect 15044 18566 15110 18582
rect 15044 18532 15060 18566
rect 15094 18532 15110 18566
rect 15044 18516 15110 18532
rect 15062 18494 15092 18516
rect 15062 16912 15092 16934
rect 15044 16896 15110 16912
rect 15044 16862 15060 16896
rect 15094 16862 15110 16896
rect 15044 16846 15110 16862
rect 15454 18566 15520 18582
rect 15454 18532 15470 18566
rect 15504 18532 15520 18566
rect 15454 18516 15520 18532
rect 15472 18494 15502 18516
rect 15472 16912 15502 16934
rect 15454 16896 15520 16912
rect 15454 16862 15470 16896
rect 15504 16862 15520 16896
rect 15454 16846 15520 16862
rect 14472 15976 14622 15994
rect 14472 15942 14566 15976
rect 14600 15942 14622 15976
rect 14472 15924 14622 15942
rect 14742 15976 14808 15992
rect 14742 15942 14758 15976
rect 14792 15942 14808 15976
rect 14472 15904 14502 15924
rect 14568 15904 14598 15924
rect 14664 15904 14694 15930
rect 14742 15926 14808 15942
rect 14934 15976 15000 15992
rect 14934 15942 14950 15976
rect 14984 15942 15000 15976
rect 14760 15904 14790 15926
rect 14856 15904 14886 15930
rect 14934 15926 15000 15942
rect 15126 15976 15192 15992
rect 15126 15942 15142 15976
rect 15176 15942 15192 15976
rect 14952 15904 14982 15926
rect 15048 15904 15078 15930
rect 15126 15926 15192 15942
rect 15144 15904 15174 15926
rect 13598 15536 13666 15554
rect 13598 15502 13616 15536
rect 13650 15502 13666 15536
rect 13598 15496 13666 15502
rect 13600 15486 13666 15496
rect 13618 15464 13648 15486
rect 13618 13882 13648 13904
rect 13600 13866 13666 13882
rect 13600 13832 13616 13866
rect 13650 13832 13666 13866
rect 13600 13816 13666 13832
rect 14472 13882 14502 13904
rect 14454 13866 14520 13882
rect 14568 13878 14598 13904
rect 14664 13882 14694 13904
rect 14454 13832 14470 13866
rect 14504 13832 14520 13866
rect 14454 13816 14520 13832
rect 14646 13866 14712 13882
rect 14760 13878 14790 13904
rect 14856 13882 14886 13904
rect 14646 13832 14662 13866
rect 14696 13832 14712 13866
rect 14646 13816 14712 13832
rect 14838 13866 14904 13882
rect 14952 13878 14982 13904
rect 15048 13882 15078 13904
rect 15144 13882 15174 13904
rect 14838 13832 14854 13866
rect 14888 13832 14904 13866
rect 14838 13816 14904 13832
rect 15030 13866 15174 13882
rect 15030 13832 15046 13866
rect 15080 13832 15174 13866
rect 15030 13816 15174 13832
rect 17142 16024 17364 16040
rect 17142 15990 17236 16024
rect 17270 15990 17364 16024
rect 17142 15969 17364 15990
rect 17142 15943 17172 15969
rect 17238 15943 17268 15969
rect 17334 15943 17364 15969
rect 17142 13917 17172 13943
rect 17238 13917 17268 13943
rect 17334 13917 17364 13943
rect 17124 13896 17382 13917
rect 17124 13862 17140 13896
rect 17174 13862 17332 13896
rect 17366 13862 17382 13896
rect 17124 13846 17382 13862
rect 17000 13310 17118 13334
rect 17000 13276 17040 13310
rect 17074 13276 17118 13310
rect 17000 13254 17118 13276
rect 13480 13181 13571 13215
rect 13480 13147 13509 13181
rect 13543 13175 13571 13181
rect 13543 13147 13598 13175
rect 13675 13172 13750 13195
rect 13480 13096 13598 13147
rect 13480 13070 13510 13096
rect 13568 13070 13598 13096
rect 13656 13171 13774 13172
rect 13656 13137 13695 13171
rect 13729 13137 13774 13171
rect 14029 13170 14104 13191
rect 14382 13172 14457 13189
rect 14735 13172 14810 13190
rect 15086 13172 15161 13190
rect 15440 13172 15515 13191
rect 15790 13173 15865 13190
rect 13656 13115 13774 13137
rect 13656 13070 13686 13115
rect 13744 13070 13774 13115
rect 14008 13167 14126 13170
rect 14008 13133 14049 13167
rect 14083 13133 14126 13167
rect 14008 13111 14126 13133
rect 13832 13070 13862 13096
rect 13920 13070 13950 13096
rect 14008 13070 14038 13111
rect 14096 13070 14126 13111
rect 14360 13165 14478 13172
rect 14360 13131 14402 13165
rect 14436 13131 14478 13165
rect 14360 13109 14478 13131
rect 14184 13070 14214 13096
rect 14272 13070 14302 13096
rect 14360 13070 14390 13109
rect 14448 13070 14478 13109
rect 14712 13166 14830 13172
rect 14712 13132 14755 13166
rect 14789 13132 14830 13166
rect 14712 13110 14830 13132
rect 14536 13070 14566 13096
rect 14624 13070 14654 13096
rect 14712 13070 14742 13110
rect 14800 13070 14830 13110
rect 15064 13166 15182 13172
rect 15064 13132 15106 13166
rect 15140 13132 15182 13166
rect 15064 13110 15182 13132
rect 14888 13070 14918 13096
rect 14976 13070 15006 13096
rect 15064 13070 15094 13110
rect 15152 13070 15182 13110
rect 15416 13167 15534 13172
rect 15416 13133 15460 13167
rect 15494 13133 15534 13167
rect 15416 13111 15534 13133
rect 15240 13070 15270 13096
rect 15328 13070 15358 13096
rect 15416 13070 15446 13111
rect 15504 13070 15534 13111
rect 15768 13166 15886 13173
rect 16142 13172 16217 13189
rect 16495 13172 16570 13189
rect 16844 13172 16919 13189
rect 15768 13132 15810 13166
rect 15844 13132 15886 13166
rect 15768 13110 15886 13132
rect 15592 13070 15622 13096
rect 15680 13070 15710 13096
rect 15768 13070 15798 13110
rect 15856 13070 15886 13110
rect 16120 13165 16238 13172
rect 16120 13131 16162 13165
rect 16196 13131 16238 13165
rect 16120 13109 16238 13131
rect 15944 13070 15974 13096
rect 16032 13070 16062 13096
rect 16120 13070 16150 13109
rect 16208 13070 16238 13109
rect 16472 13165 16590 13172
rect 16472 13131 16515 13165
rect 16549 13131 16590 13165
rect 16472 13109 16590 13131
rect 16296 13070 16326 13096
rect 16384 13070 16414 13096
rect 16472 13070 16502 13109
rect 16560 13070 16590 13109
rect 16824 13165 16942 13172
rect 16824 13131 16864 13165
rect 16898 13131 16942 13165
rect 16824 13109 16942 13131
rect 16648 13070 16678 13096
rect 16736 13070 16766 13096
rect 16824 13070 16854 13109
rect 16912 13070 16942 13109
rect 17000 13070 17030 13254
rect 17088 13070 17118 13254
rect 17198 13173 17273 13189
rect 17176 13165 17294 13173
rect 17176 13131 17218 13165
rect 17252 13131 17294 13165
rect 17371 13165 17446 13189
rect 17371 13164 17391 13165
rect 17176 13109 17294 13131
rect 17176 13070 17206 13109
rect 17264 13070 17294 13109
rect 17352 13131 17391 13164
rect 17425 13164 17446 13165
rect 17425 13131 17470 13164
rect 17352 13109 17470 13131
rect 17352 13070 17382 13109
rect 17440 13070 17470 13109
rect 13480 11020 13510 11070
rect 13568 11020 13598 11070
rect 13656 11044 13686 11070
rect 13744 11044 13774 11070
rect 13480 10996 13598 11020
rect 13480 10970 13517 10996
rect 13497 10962 13517 10970
rect 13551 10970 13598 10996
rect 13832 11014 13862 11070
rect 13920 11014 13950 11070
rect 14008 11044 14038 11070
rect 14096 11044 14126 11070
rect 13832 10990 13950 11014
rect 13551 10962 13572 10970
rect 13832 10969 13867 10990
rect 13497 10940 13572 10962
rect 13847 10956 13867 10969
rect 13901 10969 13950 10990
rect 14184 11017 14214 11070
rect 14272 11017 14302 11070
rect 14360 11044 14390 11070
rect 14448 11044 14478 11070
rect 14184 10993 14302 11017
rect 14184 10969 14225 10993
rect 13901 10956 13922 10969
rect 13847 10934 13922 10956
rect 14205 10959 14225 10969
rect 14259 10969 14302 10993
rect 14536 11017 14566 11070
rect 14624 11017 14654 11070
rect 14712 11044 14742 11070
rect 14800 11044 14830 11070
rect 14536 10993 14654 11017
rect 14536 10969 14573 10993
rect 14259 10959 14280 10969
rect 14205 10937 14280 10959
rect 14553 10959 14573 10969
rect 14607 10969 14654 10993
rect 14888 11017 14918 11070
rect 14976 11017 15006 11070
rect 15064 11044 15094 11070
rect 15152 11044 15182 11070
rect 14888 10993 15006 11017
rect 14888 10970 14924 10993
rect 14607 10959 14628 10969
rect 14553 10937 14628 10959
rect 14904 10959 14924 10970
rect 14958 10970 15006 10993
rect 15240 11016 15270 11070
rect 15328 11016 15358 11070
rect 15416 11044 15446 11070
rect 15504 11044 15534 11070
rect 15240 10992 15358 11016
rect 15240 10970 15275 10992
rect 14958 10959 14979 10970
rect 14904 10937 14979 10959
rect 15255 10958 15275 10970
rect 15309 10970 15358 10992
rect 15592 11014 15622 11070
rect 15680 11014 15710 11070
rect 15768 11044 15798 11070
rect 15856 11044 15886 11070
rect 15592 10990 15710 11014
rect 15592 10971 15626 10990
rect 15309 10958 15330 10970
rect 15255 10936 15330 10958
rect 15606 10956 15626 10971
rect 15660 10971 15710 10990
rect 15944 11017 15974 11070
rect 16032 11017 16062 11070
rect 16120 11044 16150 11070
rect 16208 11044 16238 11070
rect 15944 10993 16062 11017
rect 15944 10971 15981 10993
rect 15660 10956 15681 10971
rect 15606 10934 15681 10956
rect 15961 10959 15981 10971
rect 16015 10971 16062 10993
rect 16296 11013 16326 11070
rect 16384 11013 16414 11070
rect 16472 11044 16502 11070
rect 16560 11044 16590 11070
rect 16296 10989 16414 11013
rect 16296 10971 16331 10989
rect 16015 10959 16036 10971
rect 15961 10937 16036 10959
rect 16311 10955 16331 10971
rect 16365 10971 16414 10989
rect 16648 11015 16678 11070
rect 16736 11015 16766 11070
rect 16824 11044 16854 11070
rect 16912 11044 16942 11070
rect 16648 10991 16766 11015
rect 16365 10955 16386 10971
rect 16648 10970 16685 10991
rect 16311 10933 16386 10955
rect 16665 10957 16685 10970
rect 16719 10970 16766 10991
rect 17000 11013 17030 11070
rect 17088 11013 17118 11070
rect 17176 11044 17206 11070
rect 17264 11044 17294 11070
rect 17000 10989 17118 11013
rect 17000 10971 17035 10989
rect 16719 10957 16740 10970
rect 16665 10935 16740 10957
rect 17015 10955 17035 10971
rect 17069 10971 17118 10989
rect 17352 11024 17382 11070
rect 17440 11024 17470 11070
rect 17352 10971 17472 11024
rect 17069 10955 17090 10971
rect 17015 10933 17090 10955
rect 17352 10937 17395 10971
rect 17429 10937 17472 10971
rect 17352 10884 17472 10937
<< polycont >>
rect 16806 24078 16840 24112
rect 16998 24078 17032 24112
rect 17190 24078 17224 24112
rect 17382 24078 17416 24112
rect 17574 24078 17608 24112
rect 14114 23188 14148 23222
rect 14306 23188 14340 23222
rect 14498 23188 14532 23222
rect 14690 23188 14724 23222
rect 14018 21078 14052 21112
rect 14210 21078 14244 21112
rect 14402 21078 14436 21112
rect 14594 21078 14628 21112
rect 15974 23236 16008 23270
rect 16710 21968 16744 22002
rect 16902 21968 16936 22002
rect 17094 21968 17128 22002
rect 17286 21968 17320 22002
rect 17478 21968 17512 22002
rect 15878 21108 15912 21142
rect 16070 21108 16104 21142
rect 14974 20484 15008 20518
rect 15166 20484 15200 20518
rect 15358 20484 15392 20518
rect 14878 19088 14912 19122
rect 15070 19088 15104 19122
rect 15262 19088 15296 19122
rect 15454 19088 15488 19122
rect 16134 19998 16168 20032
rect 16038 19088 16072 19122
rect 16230 19088 16264 19122
rect 15060 18532 15094 18566
rect 15060 16862 15094 16896
rect 15470 18532 15504 18566
rect 15470 16862 15504 16896
rect 14566 15942 14600 15976
rect 14758 15942 14792 15976
rect 14950 15942 14984 15976
rect 15142 15942 15176 15976
rect 13616 15502 13650 15536
rect 13616 13832 13650 13866
rect 14470 13832 14504 13866
rect 14662 13832 14696 13866
rect 14854 13832 14888 13866
rect 15046 13832 15080 13866
rect 17236 15990 17270 16024
rect 17140 13862 17174 13896
rect 17332 13862 17366 13896
rect 17040 13276 17074 13310
rect 13509 13147 13543 13181
rect 13695 13137 13729 13171
rect 14049 13133 14083 13167
rect 14402 13131 14436 13165
rect 14755 13132 14789 13166
rect 15106 13132 15140 13166
rect 15460 13133 15494 13167
rect 15810 13132 15844 13166
rect 16162 13131 16196 13165
rect 16515 13131 16549 13165
rect 16864 13131 16898 13165
rect 17218 13131 17252 13165
rect 17391 13131 17425 13165
rect 13517 10962 13551 10996
rect 13867 10956 13901 10990
rect 14225 10959 14259 10993
rect 14573 10959 14607 10993
rect 14924 10959 14958 10993
rect 15275 10958 15309 10992
rect 15626 10956 15660 10990
rect 15981 10959 16015 10993
rect 16331 10955 16365 10989
rect 16685 10957 16719 10991
rect 17035 10955 17069 10989
rect 17395 10937 17429 10971
<< xpolycontact >>
rect 13046 24546 13478 24616
rect 16478 24546 16910 24616
rect 13076 23866 13508 23936
rect 14308 23866 14740 23936
rect 13486 21638 13556 22070
rect 13486 21106 13556 21538
rect 15306 22798 15376 23230
rect 15306 21126 15376 21558
rect 13312 19592 13744 19730
rect 13882 19592 14314 19730
rect 13312 19206 13744 19344
rect 13882 19206 14314 19344
rect 13312 18820 13744 18958
rect 13882 18820 14314 18958
rect 16786 20918 16856 21350
rect 16786 18886 16856 19318
rect 13312 18434 13744 18572
rect 13882 18434 14314 18572
rect 13312 18048 13744 18186
rect 13882 18048 14314 18186
rect 13312 17662 13744 17800
rect 13882 17662 14314 17800
rect 13312 17276 13744 17414
rect 13882 17276 14314 17414
rect 13312 16890 13744 17028
rect 13882 16890 14314 17028
rect 14642 17422 14712 17854
rect 14642 16890 14712 17322
rect 15862 17422 15932 17854
rect 15862 16890 15932 17322
rect 16254 18123 16324 18555
rect 16254 16891 16324 17323
rect 17396 20938 17466 21370
rect 17396 17506 17466 17938
rect 16148 15532 16218 15964
rect 16148 13860 16218 14292
<< ppolyres >>
rect 13478 24546 16478 24616
rect 13508 23866 14308 23936
rect 13486 21538 13556 21638
rect 15306 21558 15376 22798
rect 13744 19592 13882 19730
rect 13744 19206 13882 19344
rect 13744 18820 13882 18958
rect 16786 19318 16856 20918
rect 13744 18434 13882 18572
rect 13744 18048 13882 18186
rect 13744 17662 13882 17800
rect 13744 17276 13882 17414
rect 13744 16890 13882 17028
rect 14642 17322 14712 17422
rect 15862 17322 15932 17422
rect 16254 17323 16324 18123
rect 17396 17938 17466 20938
rect 16148 14292 16218 15532
<< ndiode >>
rect 16788 18330 16878 18358
rect 16788 18296 16816 18330
rect 16850 18296 16878 18330
rect 16788 18268 16878 18296
<< ndiodec >>
rect 16816 18296 16850 18330
<< locali >>
rect 14004 28815 16526 28932
rect 14004 27701 14128 28815
rect 16394 27701 16526 28815
rect 14004 25334 16526 27701
rect 12670 24852 17790 25334
rect 12670 23542 12834 24852
rect 13049 24746 13484 24749
rect 12916 24712 13023 24746
rect 13057 24712 13091 24746
rect 13125 24712 13159 24746
rect 13193 24712 13227 24746
rect 13261 24712 13295 24746
rect 13329 24712 13363 24746
rect 13397 24712 13431 24746
rect 13465 24712 13499 24746
rect 13533 24712 13567 24746
rect 13601 24712 13635 24746
rect 13669 24712 13703 24746
rect 13737 24712 13771 24746
rect 13805 24712 13839 24746
rect 13873 24712 13907 24746
rect 13941 24712 13975 24746
rect 14009 24712 14043 24746
rect 14077 24712 14111 24746
rect 14145 24712 14179 24746
rect 14213 24712 14247 24746
rect 14281 24712 14315 24746
rect 14349 24712 14383 24746
rect 14417 24712 14451 24746
rect 14485 24712 14519 24746
rect 14553 24712 14587 24746
rect 14621 24712 14655 24746
rect 14689 24712 14723 24746
rect 14757 24712 14791 24746
rect 14825 24712 14859 24746
rect 14893 24712 14927 24746
rect 14961 24712 14995 24746
rect 15029 24712 15063 24746
rect 15097 24712 15131 24746
rect 15165 24712 15199 24746
rect 15233 24712 15267 24746
rect 15301 24712 15335 24746
rect 15369 24712 15403 24746
rect 15437 24712 15471 24746
rect 15505 24712 15539 24746
rect 15573 24712 15607 24746
rect 15641 24712 15675 24746
rect 15709 24712 15743 24746
rect 15777 24712 15811 24746
rect 15845 24712 15879 24746
rect 15913 24712 15947 24746
rect 15981 24712 16015 24746
rect 16049 24712 16083 24746
rect 16117 24712 16151 24746
rect 16185 24712 16219 24746
rect 16253 24712 16287 24746
rect 16321 24712 16355 24746
rect 16389 24712 16423 24746
rect 16457 24712 16491 24746
rect 16525 24712 16559 24746
rect 16593 24712 16627 24746
rect 16661 24712 16695 24746
rect 16729 24712 16763 24746
rect 16797 24712 16831 24746
rect 16865 24712 16899 24746
rect 16933 24712 17040 24746
rect 12916 24632 12950 24712
rect 13049 24616 13484 24712
rect 17006 24632 17040 24712
rect 12916 24564 12950 24598
rect 13478 24546 13484 24616
rect 17006 24564 17040 24598
rect 13049 24541 13484 24546
rect 12916 24450 12950 24530
rect 17006 24450 17040 24530
rect 12916 24416 13023 24450
rect 13057 24416 13091 24450
rect 13125 24416 13159 24450
rect 13193 24416 13227 24450
rect 13261 24416 13295 24450
rect 13329 24416 13363 24450
rect 13397 24416 13431 24450
rect 13465 24416 13499 24450
rect 13533 24416 13567 24450
rect 13601 24416 13635 24450
rect 13669 24416 13703 24450
rect 13737 24416 13771 24450
rect 13805 24416 13839 24450
rect 13873 24416 13907 24450
rect 13941 24416 13975 24450
rect 14009 24416 14043 24450
rect 14077 24416 14111 24450
rect 14145 24416 14179 24450
rect 14213 24416 14247 24450
rect 14281 24416 14315 24450
rect 14349 24416 14383 24450
rect 14417 24416 14451 24450
rect 14485 24416 14519 24450
rect 14553 24416 14587 24450
rect 14621 24416 14655 24450
rect 14689 24416 14723 24450
rect 14757 24416 14791 24450
rect 14825 24416 14859 24450
rect 14893 24416 14927 24450
rect 14961 24416 14995 24450
rect 15029 24416 15063 24450
rect 15097 24416 15131 24450
rect 15165 24416 15199 24450
rect 15233 24416 15267 24450
rect 15301 24416 15335 24450
rect 15369 24416 15403 24450
rect 15437 24416 15471 24450
rect 15505 24416 15539 24450
rect 15573 24416 15607 24450
rect 15641 24416 15675 24450
rect 15709 24416 15743 24450
rect 15777 24416 15811 24450
rect 15845 24416 15879 24450
rect 15913 24416 15947 24450
rect 15981 24416 16015 24450
rect 16049 24416 16083 24450
rect 16117 24416 16151 24450
rect 16185 24416 16219 24450
rect 16253 24416 16287 24450
rect 16321 24416 16355 24450
rect 16389 24416 16423 24450
rect 16457 24416 16491 24450
rect 16525 24416 16559 24450
rect 16593 24416 16627 24450
rect 16661 24416 16695 24450
rect 16729 24416 16763 24450
rect 16797 24416 16831 24450
rect 16865 24416 16899 24450
rect 16933 24416 17040 24450
rect 16548 24180 16666 24214
rect 16700 24180 16734 24214
rect 16768 24180 16802 24214
rect 16836 24180 16870 24214
rect 16904 24180 16938 24214
rect 16972 24180 17006 24214
rect 17040 24180 17074 24214
rect 17108 24180 17142 24214
rect 17176 24180 17210 24214
rect 17244 24180 17278 24214
rect 17312 24180 17346 24214
rect 17380 24180 17414 24214
rect 17448 24180 17482 24214
rect 17516 24180 17550 24214
rect 17584 24180 17618 24214
rect 17652 24180 17770 24214
rect 16548 24111 16582 24180
rect 16790 24078 16806 24112
rect 16840 24078 16856 24112
rect 16982 24078 16998 24112
rect 17032 24078 17048 24112
rect 17174 24078 17190 24112
rect 17224 24078 17240 24112
rect 17366 24078 17382 24112
rect 17416 24078 17432 24112
rect 17558 24078 17574 24112
rect 17608 24078 17624 24112
rect 17736 24111 17770 24180
rect 12946 24032 13075 24066
rect 13109 24032 13143 24066
rect 13177 24032 13211 24066
rect 13245 24032 13279 24066
rect 13313 24032 13347 24066
rect 13381 24032 13415 24066
rect 13449 24032 13483 24066
rect 13517 24032 13551 24066
rect 13585 24032 13619 24066
rect 13653 24032 13687 24066
rect 13721 24032 13755 24066
rect 13789 24032 13823 24066
rect 13857 24032 13891 24066
rect 13925 24032 13959 24066
rect 13993 24032 14027 24066
rect 14061 24032 14095 24066
rect 14129 24032 14163 24066
rect 14197 24032 14231 24066
rect 14265 24032 14299 24066
rect 14333 24032 14367 24066
rect 14401 24032 14435 24066
rect 14469 24032 14503 24066
rect 14537 24032 14571 24066
rect 14605 24032 14639 24066
rect 14673 24032 14707 24066
rect 14741 24032 14870 24066
rect 12946 23952 12980 24032
rect 14836 23952 14870 24032
rect 12946 23884 12980 23918
rect 14836 23884 14870 23918
rect 12946 23770 12980 23850
rect 14836 23770 14870 23850
rect 12946 23736 13075 23770
rect 13109 23736 13143 23770
rect 13177 23736 13211 23770
rect 13245 23736 13279 23770
rect 13313 23736 13347 23770
rect 13381 23736 13415 23770
rect 13449 23736 13483 23770
rect 13517 23736 13551 23770
rect 13585 23736 13619 23770
rect 13653 23736 13687 23770
rect 13721 23736 13755 23770
rect 13789 23736 13823 23770
rect 13857 23736 13891 23770
rect 13925 23736 13959 23770
rect 13993 23736 14027 23770
rect 14061 23736 14095 23770
rect 14129 23736 14163 23770
rect 14197 23736 14231 23770
rect 14265 23736 14299 23770
rect 14333 23736 14367 23770
rect 14401 23736 14435 23770
rect 14469 23736 14503 23770
rect 14537 23736 14571 23770
rect 14605 23736 14639 23770
rect 14673 23736 14707 23770
rect 14741 23736 14870 23770
rect 16548 24043 16582 24077
rect 16548 23975 16582 24009
rect 16548 23907 16582 23941
rect 16548 23839 16582 23873
rect 16548 23771 16582 23805
rect 16548 23703 16582 23737
rect 16548 23635 16582 23669
rect 13300 23580 15938 23584
rect 12926 23579 15938 23580
rect 16270 23579 16450 23580
rect 12926 23548 16450 23579
rect 12926 23542 16307 23548
rect 12670 23523 16307 23542
rect 12670 23417 13111 23523
rect 13289 23442 16307 23523
rect 16413 23442 16450 23548
rect 13289 23417 16450 23442
rect 12670 23414 16450 23417
rect 12670 23378 13310 23414
rect 12926 23372 13310 23378
rect 15709 23410 16450 23414
rect 16548 23567 16582 23601
rect 16548 23499 16582 23533
rect 16548 23431 16582 23465
rect 15709 23372 16448 23410
rect 15176 23326 15290 23360
rect 15324 23326 15358 23360
rect 15392 23326 15506 23360
rect 15709 23338 15838 23372
rect 15872 23338 15906 23372
rect 15940 23338 15974 23372
rect 16008 23338 16042 23372
rect 16076 23338 16110 23372
rect 16144 23338 16448 23372
rect 15709 23332 16448 23338
rect 16548 23363 16582 23397
rect 13856 23290 13980 23324
rect 14014 23290 14048 23324
rect 14082 23290 14116 23324
rect 14150 23290 14184 23324
rect 14218 23290 14252 23324
rect 14286 23290 14320 23324
rect 14354 23290 14388 23324
rect 14422 23290 14456 23324
rect 14490 23290 14524 23324
rect 14558 23290 14592 23324
rect 14626 23290 14660 23324
rect 14694 23290 14728 23324
rect 14762 23290 14886 23324
rect 13856 23221 13890 23290
rect 14098 23188 14114 23222
rect 14148 23188 14164 23222
rect 14290 23188 14306 23222
rect 14340 23188 14356 23222
rect 14482 23188 14498 23222
rect 14532 23188 14548 23222
rect 14674 23188 14690 23222
rect 14724 23188 14740 23222
rect 14852 23221 14886 23290
rect 13856 23153 13890 23187
rect 13856 23085 13890 23119
rect 13856 23017 13890 23051
rect 13856 22949 13890 22983
rect 13856 22881 13890 22915
rect 13856 22813 13890 22847
rect 13856 22745 13890 22779
rect 13856 22677 13890 22711
rect 13856 22609 13890 22643
rect 13856 22541 13890 22575
rect 13856 22473 13890 22507
rect 13856 22405 13890 22439
rect 13856 22337 13890 22371
rect 13856 22269 13890 22303
rect 13856 22201 13890 22235
rect 13356 22166 13470 22200
rect 13504 22166 13538 22200
rect 13572 22166 13686 22200
rect 13356 22081 13390 22166
rect 13652 22081 13686 22166
rect 13356 22013 13390 22047
rect 13356 21945 13390 21979
rect 13356 21877 13390 21911
rect 13356 21809 13390 21843
rect 13356 21741 13390 21775
rect 13356 21673 13390 21707
rect 13356 21605 13390 21639
rect 13652 22013 13686 22047
rect 13652 21945 13686 21979
rect 13652 21877 13686 21911
rect 13652 21809 13686 21843
rect 13652 21741 13686 21775
rect 13652 21673 13686 21707
rect 13356 21537 13390 21571
rect 13652 21605 13686 21639
rect 13356 21469 13390 21503
rect 13356 21401 13390 21435
rect 13356 21333 13390 21367
rect 13356 21265 13390 21299
rect 13356 21197 13390 21231
rect 13356 21129 13390 21163
rect 13652 21537 13686 21571
rect 13652 21469 13686 21503
rect 13652 21401 13686 21435
rect 13652 21333 13686 21367
rect 13652 21265 13686 21299
rect 13652 21197 13686 21231
rect 13652 21129 13686 21163
rect 13356 21010 13390 21095
rect 13652 21010 13686 21095
rect 13356 20976 13470 21010
rect 13504 20976 13538 21010
rect 13572 20976 13686 21010
rect 13856 22133 13890 22167
rect 13856 22065 13890 22099
rect 13856 21997 13890 22031
rect 13856 21929 13890 21963
rect 13856 21861 13890 21895
rect 13856 21793 13890 21827
rect 13856 21725 13890 21759
rect 13856 21657 13890 21691
rect 13856 21589 13890 21623
rect 13856 21521 13890 21555
rect 13856 21453 13890 21487
rect 13856 21385 13890 21419
rect 13856 21317 13890 21351
rect 13856 21249 13890 21283
rect 13856 21181 13890 21215
rect 13856 21113 13890 21147
rect 13970 23119 14004 23154
rect 13970 23051 14004 23069
rect 13970 22983 14004 22997
rect 13970 22915 14004 22925
rect 13970 22847 14004 22853
rect 13970 22779 14004 22781
rect 13970 22743 14004 22745
rect 13970 22671 14004 22677
rect 13970 22599 14004 22609
rect 13970 22527 14004 22541
rect 13970 22455 14004 22473
rect 13970 22383 14004 22405
rect 13970 22311 14004 22337
rect 13970 22239 14004 22269
rect 13970 22167 14004 22201
rect 13970 22099 14004 22133
rect 13970 22031 14004 22061
rect 13970 21963 14004 21989
rect 13970 21895 14004 21917
rect 13970 21827 14004 21845
rect 13970 21759 14004 21773
rect 13970 21691 14004 21701
rect 13970 21623 14004 21629
rect 13970 21555 14004 21557
rect 13970 21519 14004 21521
rect 13970 21447 14004 21453
rect 13970 21375 14004 21385
rect 13970 21303 14004 21317
rect 13970 21231 14004 21249
rect 13970 21146 14004 21181
rect 14066 23119 14100 23154
rect 14066 23051 14100 23069
rect 14066 22983 14100 22997
rect 14066 22915 14100 22925
rect 14066 22847 14100 22853
rect 14066 22779 14100 22781
rect 14066 22743 14100 22745
rect 14066 22671 14100 22677
rect 14066 22599 14100 22609
rect 14066 22527 14100 22541
rect 14066 22455 14100 22473
rect 14066 22383 14100 22405
rect 14066 22311 14100 22337
rect 14066 22239 14100 22269
rect 14066 22167 14100 22201
rect 14066 22099 14100 22133
rect 14066 22031 14100 22061
rect 14066 21963 14100 21989
rect 14066 21895 14100 21917
rect 14066 21827 14100 21845
rect 14066 21759 14100 21773
rect 14066 21691 14100 21701
rect 14066 21623 14100 21629
rect 14066 21555 14100 21557
rect 14066 21519 14100 21521
rect 14066 21447 14100 21453
rect 14066 21375 14100 21385
rect 14066 21303 14100 21317
rect 14066 21231 14100 21249
rect 14066 21146 14100 21181
rect 14162 23119 14196 23154
rect 14162 23051 14196 23069
rect 14162 22983 14196 22997
rect 14162 22915 14196 22925
rect 14162 22847 14196 22853
rect 14162 22779 14196 22781
rect 14162 22743 14196 22745
rect 14162 22671 14196 22677
rect 14162 22599 14196 22609
rect 14162 22527 14196 22541
rect 14162 22455 14196 22473
rect 14162 22383 14196 22405
rect 14162 22311 14196 22337
rect 14162 22239 14196 22269
rect 14162 22167 14196 22201
rect 14162 22099 14196 22133
rect 14162 22031 14196 22061
rect 14162 21963 14196 21989
rect 14162 21895 14196 21917
rect 14162 21827 14196 21845
rect 14162 21759 14196 21773
rect 14162 21691 14196 21701
rect 14162 21623 14196 21629
rect 14162 21555 14196 21557
rect 14162 21519 14196 21521
rect 14162 21447 14196 21453
rect 14162 21375 14196 21385
rect 14162 21303 14196 21317
rect 14162 21231 14196 21249
rect 14162 21146 14196 21181
rect 14258 23119 14292 23154
rect 14258 23051 14292 23069
rect 14258 22983 14292 22997
rect 14258 22915 14292 22925
rect 14258 22847 14292 22853
rect 14258 22779 14292 22781
rect 14258 22743 14292 22745
rect 14258 22671 14292 22677
rect 14258 22599 14292 22609
rect 14258 22527 14292 22541
rect 14258 22455 14292 22473
rect 14258 22383 14292 22405
rect 14258 22311 14292 22337
rect 14258 22239 14292 22269
rect 14258 22167 14292 22201
rect 14258 22099 14292 22133
rect 14258 22031 14292 22061
rect 14258 21963 14292 21989
rect 14258 21895 14292 21917
rect 14258 21827 14292 21845
rect 14258 21759 14292 21773
rect 14258 21691 14292 21701
rect 14258 21623 14292 21629
rect 14258 21555 14292 21557
rect 14258 21519 14292 21521
rect 14258 21447 14292 21453
rect 14258 21375 14292 21385
rect 14258 21303 14292 21317
rect 14258 21231 14292 21249
rect 14258 21146 14292 21181
rect 14354 23119 14388 23154
rect 14354 23051 14388 23069
rect 14354 22983 14388 22997
rect 14354 22915 14388 22925
rect 14354 22847 14388 22853
rect 14354 22779 14388 22781
rect 14354 22743 14388 22745
rect 14354 22671 14388 22677
rect 14354 22599 14388 22609
rect 14354 22527 14388 22541
rect 14354 22455 14388 22473
rect 14354 22383 14388 22405
rect 14354 22311 14388 22337
rect 14354 22239 14388 22269
rect 14354 22167 14388 22201
rect 14354 22099 14388 22133
rect 14354 22031 14388 22061
rect 14354 21963 14388 21989
rect 14354 21895 14388 21917
rect 14354 21827 14388 21845
rect 14354 21759 14388 21773
rect 14354 21691 14388 21701
rect 14354 21623 14388 21629
rect 14354 21555 14388 21557
rect 14354 21519 14388 21521
rect 14354 21447 14388 21453
rect 14354 21375 14388 21385
rect 14354 21303 14388 21317
rect 14354 21231 14388 21249
rect 14354 21146 14388 21181
rect 14450 23119 14484 23154
rect 14450 23051 14484 23069
rect 14450 22983 14484 22997
rect 14450 22915 14484 22925
rect 14450 22847 14484 22853
rect 14450 22779 14484 22781
rect 14450 22743 14484 22745
rect 14450 22671 14484 22677
rect 14450 22599 14484 22609
rect 14450 22527 14484 22541
rect 14450 22455 14484 22473
rect 14450 22383 14484 22405
rect 14450 22311 14484 22337
rect 14450 22239 14484 22269
rect 14450 22167 14484 22201
rect 14450 22099 14484 22133
rect 14450 22031 14484 22061
rect 14450 21963 14484 21989
rect 14450 21895 14484 21917
rect 14450 21827 14484 21845
rect 14450 21759 14484 21773
rect 14450 21691 14484 21701
rect 14450 21623 14484 21629
rect 14450 21555 14484 21557
rect 14450 21519 14484 21521
rect 14450 21447 14484 21453
rect 14450 21375 14484 21385
rect 14450 21303 14484 21317
rect 14450 21231 14484 21249
rect 14450 21146 14484 21181
rect 14546 23119 14580 23154
rect 14546 23051 14580 23069
rect 14546 22983 14580 22997
rect 14546 22915 14580 22925
rect 14546 22847 14580 22853
rect 14546 22779 14580 22781
rect 14546 22743 14580 22745
rect 14546 22671 14580 22677
rect 14546 22599 14580 22609
rect 14546 22527 14580 22541
rect 14546 22455 14580 22473
rect 14546 22383 14580 22405
rect 14546 22311 14580 22337
rect 14546 22239 14580 22269
rect 14546 22167 14580 22201
rect 14546 22099 14580 22133
rect 14546 22031 14580 22061
rect 14546 21963 14580 21989
rect 14546 21895 14580 21917
rect 14546 21827 14580 21845
rect 14546 21759 14580 21773
rect 14546 21691 14580 21701
rect 14546 21623 14580 21629
rect 14546 21555 14580 21557
rect 14546 21519 14580 21521
rect 14546 21447 14580 21453
rect 14546 21375 14580 21385
rect 14546 21303 14580 21317
rect 14546 21231 14580 21249
rect 14546 21146 14580 21181
rect 14642 23119 14676 23154
rect 14642 23051 14676 23069
rect 14642 22983 14676 22997
rect 14642 22915 14676 22925
rect 14642 22847 14676 22853
rect 14642 22779 14676 22781
rect 14642 22743 14676 22745
rect 14642 22671 14676 22677
rect 14642 22599 14676 22609
rect 14642 22527 14676 22541
rect 14642 22455 14676 22473
rect 14642 22383 14676 22405
rect 14642 22311 14676 22337
rect 14642 22239 14676 22269
rect 14642 22167 14676 22201
rect 14642 22099 14676 22133
rect 14642 22031 14676 22061
rect 14642 21963 14676 21989
rect 14642 21895 14676 21917
rect 14642 21827 14676 21845
rect 14642 21759 14676 21773
rect 14642 21691 14676 21701
rect 14642 21623 14676 21629
rect 14642 21555 14676 21557
rect 14642 21519 14676 21521
rect 14642 21447 14676 21453
rect 14642 21375 14676 21385
rect 14642 21303 14676 21317
rect 14642 21231 14676 21249
rect 14642 21146 14676 21181
rect 14738 23119 14772 23154
rect 14852 23153 14886 23187
rect 14738 23051 14772 23069
rect 14820 23119 14852 23150
rect 15176 23249 15210 23326
rect 15472 23249 15506 23326
rect 15176 23181 15210 23215
rect 14886 23119 14910 23150
rect 14820 23107 14910 23119
rect 14820 23073 14848 23107
rect 14882 23085 14910 23107
rect 14820 23051 14852 23073
rect 14886 23051 14910 23085
rect 14820 23030 14910 23051
rect 15176 23113 15210 23147
rect 15176 23045 15210 23079
rect 14738 22983 14772 22997
rect 14738 22915 14772 22925
rect 14738 22847 14772 22853
rect 14738 22779 14772 22781
rect 14738 22743 14772 22745
rect 14738 22671 14772 22677
rect 14738 22599 14772 22609
rect 14738 22527 14772 22541
rect 14738 22455 14772 22473
rect 14738 22383 14772 22405
rect 14738 22311 14772 22337
rect 14738 22239 14772 22269
rect 14738 22167 14772 22201
rect 14738 22099 14772 22133
rect 14738 22031 14772 22061
rect 14738 21963 14772 21989
rect 14738 21895 14772 21917
rect 14738 21827 14772 21845
rect 14738 21759 14772 21773
rect 14738 21691 14772 21701
rect 14738 21623 14772 21629
rect 14738 21555 14772 21557
rect 14738 21519 14772 21521
rect 14738 21447 14772 21453
rect 14738 21375 14772 21385
rect 14738 21303 14772 21317
rect 14738 21231 14772 21249
rect 14738 21146 14772 21181
rect 14852 23017 14886 23030
rect 14852 22949 14886 22983
rect 14852 22881 14886 22915
rect 14852 22813 14886 22847
rect 14852 22745 14886 22779
rect 14852 22677 14886 22711
rect 14852 22609 14886 22643
rect 14852 22541 14886 22575
rect 14852 22473 14886 22507
rect 14852 22405 14886 22439
rect 14852 22337 14886 22371
rect 14852 22269 14886 22303
rect 14852 22201 14886 22235
rect 14852 22133 14886 22167
rect 14852 22065 14886 22099
rect 14852 21997 14886 22031
rect 14852 21929 14886 21963
rect 14852 21861 14886 21895
rect 14852 21793 14886 21827
rect 14852 21725 14886 21759
rect 14852 21657 14886 21691
rect 14852 21589 14886 21623
rect 14852 21521 14886 21555
rect 14852 21453 14886 21487
rect 14852 21385 14886 21419
rect 14852 21317 14886 21351
rect 14852 21249 14886 21283
rect 14852 21181 14886 21215
rect 14852 21113 14886 21147
rect 13856 21010 13890 21079
rect 14002 21078 14018 21112
rect 14052 21078 14068 21112
rect 14194 21078 14210 21112
rect 14244 21078 14260 21112
rect 14386 21078 14402 21112
rect 14436 21078 14452 21112
rect 14578 21078 14594 21112
rect 14628 21078 14644 21112
rect 14852 21010 14886 21079
rect 13856 20976 13980 21010
rect 14014 20976 14048 21010
rect 14082 20976 14116 21010
rect 14150 20976 14184 21010
rect 14218 20976 14252 21010
rect 14286 20976 14320 21010
rect 14354 20976 14388 21010
rect 14422 20976 14456 21010
rect 14490 20976 14524 21010
rect 14558 20976 14592 21010
rect 14626 20976 14660 21010
rect 14694 20976 14728 21010
rect 14762 20976 14886 21010
rect 15176 22977 15210 23011
rect 15176 22909 15210 22943
rect 15176 22841 15210 22875
rect 15176 22773 15210 22807
rect 15472 23181 15506 23215
rect 15472 23113 15506 23147
rect 15472 23045 15506 23079
rect 15472 22977 15506 23011
rect 15472 22909 15506 22943
rect 15472 22841 15506 22875
rect 15176 22705 15210 22739
rect 15176 22637 15210 22671
rect 15176 22569 15210 22603
rect 15176 22501 15210 22535
rect 15176 22433 15210 22467
rect 15176 22365 15210 22399
rect 15176 22297 15210 22331
rect 15176 22229 15210 22263
rect 15176 22161 15210 22195
rect 15176 22093 15210 22127
rect 15176 22025 15210 22059
rect 15176 21957 15210 21991
rect 15176 21889 15210 21923
rect 15176 21821 15210 21855
rect 15176 21753 15210 21787
rect 15176 21685 15210 21719
rect 15176 21617 15210 21651
rect 15176 21549 15210 21583
rect 15472 22773 15506 22807
rect 15472 22705 15506 22739
rect 15472 22637 15506 22671
rect 15472 22569 15506 22603
rect 15472 22501 15506 22535
rect 15472 22433 15506 22467
rect 15472 22365 15506 22399
rect 15472 22297 15506 22331
rect 15472 22229 15506 22263
rect 15472 22161 15506 22195
rect 15472 22093 15506 22127
rect 15472 22025 15506 22059
rect 15472 21957 15506 21991
rect 15472 21889 15506 21923
rect 15472 21821 15506 21855
rect 15472 21753 15506 21787
rect 15472 21685 15506 21719
rect 15472 21617 15506 21651
rect 15176 21481 15210 21515
rect 15176 21413 15210 21447
rect 15176 21345 15210 21379
rect 15176 21277 15210 21311
rect 15176 21209 15210 21243
rect 15176 21141 15210 21175
rect 15472 21549 15506 21583
rect 15472 21481 15506 21515
rect 15472 21413 15506 21447
rect 15472 21345 15506 21379
rect 15472 21277 15506 21311
rect 15472 21209 15506 21243
rect 15472 21141 15506 21175
rect 15176 21030 15210 21107
rect 15472 21030 15506 21107
rect 15176 20996 15290 21030
rect 15324 20996 15358 21030
rect 15392 20996 15506 21030
rect 15716 23260 15750 23332
rect 15958 23236 15974 23270
rect 16008 23236 16024 23270
rect 16232 23260 16266 23332
rect 15716 23192 15750 23226
rect 15716 23124 15750 23158
rect 15716 23056 15750 23090
rect 15716 22988 15750 23022
rect 15716 22920 15750 22954
rect 15716 22852 15750 22886
rect 15716 22784 15750 22818
rect 15716 22716 15750 22750
rect 15716 22648 15750 22682
rect 15716 22580 15750 22614
rect 15716 22512 15750 22546
rect 15716 22444 15750 22478
rect 15716 22376 15750 22410
rect 15716 22308 15750 22342
rect 15716 22240 15750 22274
rect 15716 22172 15750 22206
rect 15716 22104 15750 22138
rect 15716 22036 15750 22070
rect 15716 21968 15750 22002
rect 15716 21900 15750 21934
rect 15716 21832 15750 21866
rect 15716 21764 15750 21798
rect 15716 21696 15750 21730
rect 15716 21628 15750 21662
rect 15716 21560 15750 21594
rect 15716 21492 15750 21526
rect 15716 21424 15750 21458
rect 15716 21356 15750 21390
rect 15716 21288 15750 21322
rect 15716 21220 15750 21254
rect 15716 21152 15750 21186
rect 15830 23158 15864 23193
rect 15830 23090 15864 23108
rect 15830 23022 15864 23036
rect 15830 22954 15864 22964
rect 15830 22886 15864 22892
rect 15830 22818 15864 22820
rect 15830 22782 15864 22784
rect 15830 22710 15864 22716
rect 15830 22638 15864 22648
rect 15830 22566 15864 22580
rect 15830 22494 15864 22512
rect 15830 22422 15864 22444
rect 15830 22350 15864 22376
rect 15830 22278 15864 22308
rect 15830 22206 15864 22240
rect 15830 22138 15864 22172
rect 15830 22070 15864 22100
rect 15830 22002 15864 22028
rect 15830 21934 15864 21956
rect 15830 21866 15864 21884
rect 15830 21798 15864 21812
rect 15830 21730 15864 21740
rect 15830 21662 15864 21668
rect 15830 21594 15864 21596
rect 15830 21558 15864 21560
rect 15830 21486 15864 21492
rect 15830 21414 15864 21424
rect 15830 21342 15864 21356
rect 15830 21270 15864 21288
rect 15830 21185 15864 21220
rect 15926 23158 15960 23193
rect 15926 23090 15960 23108
rect 15926 23022 15960 23036
rect 15926 22954 15960 22964
rect 15926 22886 15960 22892
rect 15926 22818 15960 22820
rect 15926 22782 15960 22784
rect 15926 22710 15960 22716
rect 15926 22638 15960 22648
rect 15926 22566 15960 22580
rect 15926 22494 15960 22512
rect 15926 22422 15960 22444
rect 15926 22350 15960 22376
rect 15926 22278 15960 22308
rect 15926 22206 15960 22240
rect 15926 22138 15960 22172
rect 15926 22070 15960 22100
rect 15926 22002 15960 22028
rect 15926 21934 15960 21956
rect 15926 21866 15960 21884
rect 15926 21798 15960 21812
rect 15926 21730 15960 21740
rect 15926 21662 15960 21668
rect 15926 21594 15960 21596
rect 15926 21558 15960 21560
rect 15926 21486 15960 21492
rect 15926 21414 15960 21424
rect 15926 21342 15960 21356
rect 15926 21270 15960 21288
rect 15926 21185 15960 21220
rect 16022 23158 16056 23193
rect 16022 23090 16056 23108
rect 16022 23022 16056 23036
rect 16022 22954 16056 22964
rect 16022 22886 16056 22892
rect 16022 22818 16056 22820
rect 16022 22782 16056 22784
rect 16022 22710 16056 22716
rect 16022 22638 16056 22648
rect 16022 22566 16056 22580
rect 16022 22494 16056 22512
rect 16022 22422 16056 22444
rect 16022 22350 16056 22376
rect 16022 22278 16056 22308
rect 16022 22206 16056 22240
rect 16022 22138 16056 22172
rect 16022 22070 16056 22100
rect 16022 22002 16056 22028
rect 16022 21934 16056 21956
rect 16022 21866 16056 21884
rect 16022 21798 16056 21812
rect 16022 21730 16056 21740
rect 16022 21662 16056 21668
rect 16022 21594 16056 21596
rect 16022 21558 16056 21560
rect 16022 21486 16056 21492
rect 16022 21414 16056 21424
rect 16022 21342 16056 21356
rect 16022 21270 16056 21288
rect 16022 21185 16056 21220
rect 16118 23190 16152 23193
rect 16232 23192 16266 23226
rect 16118 23158 16232 23190
rect 16548 23295 16582 23329
rect 16548 23227 16582 23261
rect 16266 23158 16270 23190
rect 16152 23124 16270 23158
rect 16152 23108 16232 23124
rect 16118 23090 16232 23108
rect 16266 23090 16270 23124
rect 16152 23070 16270 23090
rect 16548 23159 16582 23193
rect 16548 23091 16582 23125
rect 16118 23022 16152 23036
rect 16118 22954 16152 22964
rect 16118 22886 16152 22892
rect 16118 22818 16152 22820
rect 16118 22782 16152 22784
rect 16118 22710 16152 22716
rect 16118 22638 16152 22648
rect 16118 22566 16152 22580
rect 16118 22494 16152 22512
rect 16118 22422 16152 22444
rect 16118 22350 16152 22376
rect 16118 22278 16152 22308
rect 16118 22206 16152 22240
rect 16118 22138 16152 22172
rect 16118 22070 16152 22100
rect 16118 22002 16152 22028
rect 16118 21934 16152 21956
rect 16118 21866 16152 21884
rect 16118 21798 16152 21812
rect 16232 23056 16266 23070
rect 16232 22988 16266 23022
rect 16232 22920 16266 22954
rect 16232 22852 16266 22886
rect 16232 22784 16266 22818
rect 16232 22716 16266 22750
rect 16232 22648 16266 22682
rect 16232 22580 16266 22614
rect 16232 22512 16266 22546
rect 16232 22444 16266 22478
rect 16232 22376 16266 22410
rect 16232 22308 16266 22342
rect 16232 22240 16266 22274
rect 16232 22172 16266 22206
rect 16232 22104 16266 22138
rect 16232 22036 16266 22070
rect 16232 21968 16266 22002
rect 16232 21900 16266 21934
rect 16548 23023 16582 23057
rect 16548 22955 16582 22989
rect 16548 22887 16582 22921
rect 16548 22819 16582 22853
rect 16548 22751 16582 22785
rect 16548 22683 16582 22717
rect 16548 22615 16582 22649
rect 16548 22547 16582 22581
rect 16548 22479 16582 22513
rect 16548 22411 16582 22445
rect 16548 22343 16582 22377
rect 16548 22275 16582 22309
rect 16548 22207 16582 22241
rect 16548 22139 16582 22173
rect 16548 22071 16582 22105
rect 16548 22003 16582 22037
rect 16662 24009 16696 24044
rect 16662 23941 16696 23959
rect 16662 23873 16696 23887
rect 16662 23805 16696 23815
rect 16662 23737 16696 23743
rect 16662 23669 16696 23671
rect 16662 23633 16696 23635
rect 16662 23561 16696 23567
rect 16662 23489 16696 23499
rect 16662 23417 16696 23431
rect 16662 23345 16696 23363
rect 16662 23273 16696 23295
rect 16662 23201 16696 23227
rect 16662 23129 16696 23159
rect 16662 23057 16696 23091
rect 16662 22989 16696 23023
rect 16662 22921 16696 22951
rect 16662 22853 16696 22879
rect 16662 22785 16696 22807
rect 16662 22717 16696 22735
rect 16662 22649 16696 22663
rect 16662 22581 16696 22591
rect 16662 22513 16696 22519
rect 16662 22445 16696 22447
rect 16662 22409 16696 22411
rect 16662 22337 16696 22343
rect 16662 22265 16696 22275
rect 16662 22193 16696 22207
rect 16662 22121 16696 22139
rect 16662 22036 16696 22071
rect 16758 24009 16792 24044
rect 16758 23941 16792 23959
rect 16758 23873 16792 23887
rect 16758 23805 16792 23815
rect 16758 23737 16792 23743
rect 16758 23669 16792 23671
rect 16758 23633 16792 23635
rect 16758 23561 16792 23567
rect 16758 23489 16792 23499
rect 16758 23417 16792 23431
rect 16758 23345 16792 23363
rect 16758 23273 16792 23295
rect 16758 23201 16792 23227
rect 16758 23129 16792 23159
rect 16758 23057 16792 23091
rect 16758 22989 16792 23023
rect 16758 22921 16792 22951
rect 16758 22853 16792 22879
rect 16758 22785 16792 22807
rect 16758 22717 16792 22735
rect 16758 22649 16792 22663
rect 16758 22581 16792 22591
rect 16758 22513 16792 22519
rect 16758 22445 16792 22447
rect 16758 22409 16792 22411
rect 16758 22337 16792 22343
rect 16758 22265 16792 22275
rect 16758 22193 16792 22207
rect 16758 22121 16792 22139
rect 16758 22036 16792 22071
rect 16854 24009 16888 24044
rect 16854 23941 16888 23959
rect 16854 23873 16888 23887
rect 16854 23805 16888 23815
rect 16854 23737 16888 23743
rect 16854 23669 16888 23671
rect 16854 23633 16888 23635
rect 16854 23561 16888 23567
rect 16854 23489 16888 23499
rect 16854 23417 16888 23431
rect 16854 23345 16888 23363
rect 16854 23273 16888 23295
rect 16854 23201 16888 23227
rect 16854 23129 16888 23159
rect 16854 23057 16888 23091
rect 16854 22989 16888 23023
rect 16854 22921 16888 22951
rect 16854 22853 16888 22879
rect 16854 22785 16888 22807
rect 16854 22717 16888 22735
rect 16854 22649 16888 22663
rect 16854 22581 16888 22591
rect 16854 22513 16888 22519
rect 16854 22445 16888 22447
rect 16854 22409 16888 22411
rect 16854 22337 16888 22343
rect 16854 22265 16888 22275
rect 16854 22193 16888 22207
rect 16854 22121 16888 22139
rect 16854 22036 16888 22071
rect 16950 24009 16984 24044
rect 16950 23941 16984 23959
rect 16950 23873 16984 23887
rect 16950 23805 16984 23815
rect 16950 23737 16984 23743
rect 16950 23669 16984 23671
rect 16950 23633 16984 23635
rect 16950 23561 16984 23567
rect 16950 23489 16984 23499
rect 16950 23417 16984 23431
rect 16950 23345 16984 23363
rect 16950 23273 16984 23295
rect 16950 23201 16984 23227
rect 16950 23129 16984 23159
rect 16950 23057 16984 23091
rect 16950 22989 16984 23023
rect 16950 22921 16984 22951
rect 16950 22853 16984 22879
rect 16950 22785 16984 22807
rect 16950 22717 16984 22735
rect 16950 22649 16984 22663
rect 16950 22581 16984 22591
rect 16950 22513 16984 22519
rect 16950 22445 16984 22447
rect 16950 22409 16984 22411
rect 16950 22337 16984 22343
rect 16950 22265 16984 22275
rect 16950 22193 16984 22207
rect 16950 22121 16984 22139
rect 16950 22036 16984 22071
rect 17046 24009 17080 24044
rect 17046 23941 17080 23959
rect 17046 23873 17080 23887
rect 17046 23805 17080 23815
rect 17046 23737 17080 23743
rect 17046 23669 17080 23671
rect 17046 23633 17080 23635
rect 17046 23561 17080 23567
rect 17046 23489 17080 23499
rect 17046 23417 17080 23431
rect 17046 23345 17080 23363
rect 17046 23273 17080 23295
rect 17046 23201 17080 23227
rect 17046 23129 17080 23159
rect 17046 23057 17080 23091
rect 17046 22989 17080 23023
rect 17046 22921 17080 22951
rect 17046 22853 17080 22879
rect 17046 22785 17080 22807
rect 17046 22717 17080 22735
rect 17046 22649 17080 22663
rect 17046 22581 17080 22591
rect 17046 22513 17080 22519
rect 17046 22445 17080 22447
rect 17046 22409 17080 22411
rect 17046 22337 17080 22343
rect 17046 22265 17080 22275
rect 17046 22193 17080 22207
rect 17046 22121 17080 22139
rect 17046 22036 17080 22071
rect 17142 24009 17176 24044
rect 17142 23941 17176 23959
rect 17142 23873 17176 23887
rect 17142 23805 17176 23815
rect 17142 23737 17176 23743
rect 17142 23669 17176 23671
rect 17142 23633 17176 23635
rect 17142 23561 17176 23567
rect 17142 23489 17176 23499
rect 17142 23417 17176 23431
rect 17142 23345 17176 23363
rect 17142 23273 17176 23295
rect 17142 23201 17176 23227
rect 17142 23129 17176 23159
rect 17142 23057 17176 23091
rect 17142 22989 17176 23023
rect 17142 22921 17176 22951
rect 17142 22853 17176 22879
rect 17142 22785 17176 22807
rect 17142 22717 17176 22735
rect 17142 22649 17176 22663
rect 17142 22581 17176 22591
rect 17142 22513 17176 22519
rect 17142 22445 17176 22447
rect 17142 22409 17176 22411
rect 17142 22337 17176 22343
rect 17142 22265 17176 22275
rect 17142 22193 17176 22207
rect 17142 22121 17176 22139
rect 17142 22036 17176 22071
rect 17238 24009 17272 24044
rect 17238 23941 17272 23959
rect 17238 23873 17272 23887
rect 17238 23805 17272 23815
rect 17238 23737 17272 23743
rect 17238 23669 17272 23671
rect 17238 23633 17272 23635
rect 17238 23561 17272 23567
rect 17238 23489 17272 23499
rect 17238 23417 17272 23431
rect 17238 23345 17272 23363
rect 17238 23273 17272 23295
rect 17238 23201 17272 23227
rect 17238 23129 17272 23159
rect 17238 23057 17272 23091
rect 17238 22989 17272 23023
rect 17238 22921 17272 22951
rect 17238 22853 17272 22879
rect 17238 22785 17272 22807
rect 17238 22717 17272 22735
rect 17238 22649 17272 22663
rect 17238 22581 17272 22591
rect 17238 22513 17272 22519
rect 17238 22445 17272 22447
rect 17238 22409 17272 22411
rect 17238 22337 17272 22343
rect 17238 22265 17272 22275
rect 17238 22193 17272 22207
rect 17238 22121 17272 22139
rect 17238 22036 17272 22071
rect 17334 24009 17368 24044
rect 17334 23941 17368 23959
rect 17334 23873 17368 23887
rect 17334 23805 17368 23815
rect 17334 23737 17368 23743
rect 17334 23669 17368 23671
rect 17334 23633 17368 23635
rect 17334 23561 17368 23567
rect 17334 23489 17368 23499
rect 17334 23417 17368 23431
rect 17334 23345 17368 23363
rect 17334 23273 17368 23295
rect 17334 23201 17368 23227
rect 17334 23129 17368 23159
rect 17334 23057 17368 23091
rect 17334 22989 17368 23023
rect 17334 22921 17368 22951
rect 17334 22853 17368 22879
rect 17334 22785 17368 22807
rect 17334 22717 17368 22735
rect 17334 22649 17368 22663
rect 17334 22581 17368 22591
rect 17334 22513 17368 22519
rect 17334 22445 17368 22447
rect 17334 22409 17368 22411
rect 17334 22337 17368 22343
rect 17334 22265 17368 22275
rect 17334 22193 17368 22207
rect 17334 22121 17368 22139
rect 17334 22036 17368 22071
rect 17430 24009 17464 24044
rect 17430 23941 17464 23959
rect 17430 23873 17464 23887
rect 17430 23805 17464 23815
rect 17430 23737 17464 23743
rect 17430 23669 17464 23671
rect 17430 23633 17464 23635
rect 17430 23561 17464 23567
rect 17430 23489 17464 23499
rect 17430 23417 17464 23431
rect 17430 23345 17464 23363
rect 17430 23273 17464 23295
rect 17430 23201 17464 23227
rect 17430 23129 17464 23159
rect 17430 23057 17464 23091
rect 17430 22989 17464 23023
rect 17430 22921 17464 22951
rect 17430 22853 17464 22879
rect 17430 22785 17464 22807
rect 17430 22717 17464 22735
rect 17430 22649 17464 22663
rect 17430 22581 17464 22591
rect 17430 22513 17464 22519
rect 17430 22445 17464 22447
rect 17430 22409 17464 22411
rect 17430 22337 17464 22343
rect 17430 22265 17464 22275
rect 17430 22193 17464 22207
rect 17430 22121 17464 22139
rect 17430 22036 17464 22071
rect 17526 24009 17560 24044
rect 17526 23941 17560 23959
rect 17526 23873 17560 23887
rect 17526 23805 17560 23815
rect 17526 23737 17560 23743
rect 17526 23669 17560 23671
rect 17526 23633 17560 23635
rect 17526 23561 17560 23567
rect 17526 23489 17560 23499
rect 17526 23417 17560 23431
rect 17526 23345 17560 23363
rect 17526 23273 17560 23295
rect 17526 23201 17560 23227
rect 17526 23129 17560 23159
rect 17526 23057 17560 23091
rect 17526 22989 17560 23023
rect 17526 22921 17560 22951
rect 17526 22853 17560 22879
rect 17526 22785 17560 22807
rect 17526 22717 17560 22735
rect 17526 22649 17560 22663
rect 17526 22581 17560 22591
rect 17526 22513 17560 22519
rect 17526 22445 17560 22447
rect 17526 22409 17560 22411
rect 17526 22337 17560 22343
rect 17526 22265 17560 22275
rect 17526 22193 17560 22207
rect 17526 22121 17560 22139
rect 17526 22036 17560 22071
rect 17622 24009 17656 24044
rect 17622 23941 17656 23959
rect 17622 23873 17656 23887
rect 17622 23805 17656 23815
rect 17622 23737 17656 23743
rect 17622 23669 17656 23671
rect 17622 23633 17656 23635
rect 17622 23561 17656 23567
rect 17622 23489 17656 23499
rect 17622 23417 17656 23431
rect 17622 23345 17656 23363
rect 17622 23273 17656 23295
rect 17622 23201 17656 23227
rect 17622 23129 17656 23159
rect 17622 23057 17656 23091
rect 17622 22989 17656 23023
rect 17622 22921 17656 22951
rect 17622 22853 17656 22879
rect 17622 22785 17656 22807
rect 17622 22717 17656 22735
rect 17622 22649 17656 22663
rect 17622 22581 17656 22591
rect 17622 22513 17656 22519
rect 17622 22445 17656 22447
rect 17622 22409 17656 22411
rect 17622 22337 17656 22343
rect 17622 22265 17656 22275
rect 17622 22193 17656 22207
rect 17622 22121 17656 22139
rect 17622 22036 17656 22071
rect 17736 24043 17770 24077
rect 17736 23975 17770 24009
rect 17736 23907 17770 23941
rect 17736 23839 17770 23873
rect 17736 23771 17770 23805
rect 17736 23703 17770 23737
rect 17736 23635 17770 23669
rect 17736 23567 17770 23601
rect 17736 23499 17770 23533
rect 17736 23431 17770 23465
rect 17736 23363 17770 23397
rect 17736 23295 17770 23329
rect 17736 23227 17770 23261
rect 17736 23159 17770 23193
rect 17736 23091 17770 23125
rect 17736 23023 17770 23057
rect 17736 22955 17770 22989
rect 17736 22887 17770 22921
rect 17736 22819 17770 22853
rect 17736 22751 17770 22785
rect 17736 22683 17770 22717
rect 17736 22615 17770 22649
rect 17736 22547 17770 22581
rect 17736 22479 17770 22513
rect 17736 22411 17770 22445
rect 17736 22343 17770 22377
rect 17736 22275 17770 22309
rect 17736 22207 17770 22241
rect 17736 22139 17770 22173
rect 17736 22071 17770 22105
rect 17736 22003 17770 22037
rect 16548 21900 16582 21969
rect 16694 21968 16710 22002
rect 16744 21968 16760 22002
rect 16886 21968 16902 22002
rect 16936 21968 16952 22002
rect 17078 21968 17094 22002
rect 17128 21968 17144 22002
rect 17270 21968 17286 22002
rect 17320 21968 17336 22002
rect 17462 21968 17478 22002
rect 17512 21968 17528 22002
rect 17736 21900 17770 21969
rect 16548 21866 16666 21900
rect 16700 21866 16734 21900
rect 16768 21866 16802 21900
rect 16836 21866 16870 21900
rect 16904 21866 16938 21900
rect 16972 21866 17006 21900
rect 17040 21866 17074 21900
rect 17108 21866 17142 21900
rect 17176 21866 17210 21900
rect 17244 21866 17278 21900
rect 17312 21866 17346 21900
rect 17380 21866 17414 21900
rect 17448 21866 17482 21900
rect 17516 21866 17550 21900
rect 17584 21866 17618 21900
rect 17652 21866 17770 21900
rect 16232 21832 16266 21866
rect 16232 21775 16266 21798
rect 16118 21730 16152 21740
rect 16118 21662 16152 21668
rect 16118 21594 16152 21596
rect 16225 21764 17635 21775
rect 16225 21730 16232 21764
rect 16266 21730 17635 21764
rect 16225 21718 17635 21730
rect 16225 21696 17387 21718
rect 16225 21662 16232 21696
rect 16266 21662 17387 21696
rect 16225 21628 17387 21662
rect 16225 21594 16232 21628
rect 16266 21612 17387 21628
rect 17493 21612 17635 21718
rect 16266 21594 17635 21612
rect 16225 21565 17635 21594
rect 16118 21558 16152 21560
rect 16118 21486 16152 21492
rect 16118 21414 16152 21424
rect 16118 21342 16152 21356
rect 16118 21270 16152 21288
rect 16118 21185 16152 21220
rect 16232 21560 16266 21565
rect 16232 21492 16266 21526
rect 16232 21424 16266 21458
rect 16232 21356 16266 21390
rect 16232 21288 16266 21322
rect 16232 21220 16266 21254
rect 16232 21152 16266 21186
rect 15716 21040 15750 21118
rect 15862 21108 15878 21142
rect 15912 21108 15928 21142
rect 16054 21108 16070 21142
rect 16104 21108 16120 21142
rect 16232 21040 16266 21118
rect 15716 21006 15838 21040
rect 15872 21006 15906 21040
rect 15940 21006 15974 21040
rect 16008 21006 16042 21040
rect 16076 21006 16110 21040
rect 16144 21006 16266 21040
rect 16656 21446 16770 21480
rect 16804 21446 16838 21480
rect 16872 21446 16986 21480
rect 16656 21359 16690 21446
rect 16952 21359 16986 21446
rect 16656 21291 16690 21325
rect 16656 21223 16690 21257
rect 16656 21155 16690 21189
rect 16656 21087 16690 21121
rect 16656 21019 16690 21053
rect 16656 20951 16690 20985
rect 16952 21291 16986 21325
rect 16952 21223 16986 21257
rect 16952 21155 16986 21189
rect 16952 21087 16986 21121
rect 16952 21019 16986 21053
rect 16952 20951 16986 20985
rect 16656 20883 16690 20917
rect 16656 20815 16690 20849
rect 16656 20747 16690 20781
rect 16656 20679 16690 20713
rect 14716 20586 14826 20620
rect 14860 20586 14894 20620
rect 14928 20586 14962 20620
rect 14996 20586 15030 20620
rect 15064 20586 15098 20620
rect 15132 20586 15166 20620
rect 15200 20586 15234 20620
rect 15268 20586 15302 20620
rect 15336 20586 15370 20620
rect 15404 20586 15438 20620
rect 15472 20586 15506 20620
rect 15540 20586 15650 20620
rect 14716 20500 14750 20586
rect 14958 20484 14974 20518
rect 15008 20484 15024 20518
rect 15150 20484 15166 20518
rect 15200 20484 15216 20518
rect 15342 20484 15358 20518
rect 15392 20484 15408 20518
rect 15616 20500 15650 20586
rect 14716 20432 14750 20466
rect 14716 20364 14750 20398
rect 14716 20296 14750 20330
rect 14716 20228 14750 20262
rect 14716 20160 14750 20194
rect 14716 20092 14750 20126
rect 14716 20024 14750 20058
rect 14716 19956 14750 19990
rect 14716 19888 14750 19922
rect 13182 19826 13286 19860
rect 13320 19826 13354 19860
rect 13388 19826 13422 19860
rect 13456 19826 13490 19860
rect 13524 19826 13558 19860
rect 13592 19826 13626 19860
rect 13660 19826 13694 19860
rect 13728 19826 13762 19860
rect 13796 19826 13830 19860
rect 13864 19826 13898 19860
rect 13932 19826 13966 19860
rect 14000 19826 14034 19860
rect 14068 19826 14102 19860
rect 14136 19826 14170 19860
rect 14204 19826 14238 19860
rect 14272 19826 14306 19860
rect 14340 19826 14444 19860
rect 13182 19755 13216 19826
rect 14410 19755 14444 19826
rect 13182 19687 13216 19721
rect 13182 19619 13216 19653
rect 14410 19687 14444 19721
rect 14410 19619 14444 19653
rect 13182 19551 13216 19585
rect 13182 19483 13216 19517
rect 13182 19415 13216 19449
rect 13182 19347 13216 19381
rect 14410 19551 14444 19585
rect 14410 19483 14444 19517
rect 14410 19415 14444 19449
rect 14410 19347 14444 19381
rect 13182 19279 13216 19313
rect 13182 19211 13216 19245
rect 14410 19279 14444 19313
rect 14410 19211 14444 19245
rect 13182 19143 13216 19177
rect 13182 19075 13216 19109
rect 13182 19007 13216 19041
rect 13182 18939 13216 18973
rect 14410 19143 14444 19177
rect 14410 19075 14444 19109
rect 14410 19007 14444 19041
rect 14716 19820 14750 19854
rect 14716 19752 14750 19786
rect 14716 19684 14750 19718
rect 14716 19616 14750 19650
rect 14716 19548 14750 19582
rect 14716 19480 14750 19514
rect 14716 19412 14750 19446
rect 14716 19344 14750 19378
rect 14716 19300 14750 19310
rect 14830 20432 14864 20450
rect 14830 20364 14864 20398
rect 14830 20296 14864 20326
rect 14830 20228 14864 20254
rect 14830 20160 14864 20182
rect 14830 20092 14864 20110
rect 14830 20024 14864 20038
rect 14830 19956 14864 19966
rect 14830 19888 14864 19894
rect 14830 19820 14864 19822
rect 14830 19784 14864 19786
rect 14830 19712 14864 19718
rect 14830 19640 14864 19650
rect 14830 19568 14864 19582
rect 14830 19496 14864 19514
rect 14830 19424 14864 19446
rect 14830 19352 14864 19378
rect 14830 19300 14864 19310
rect 14926 20432 14960 20450
rect 14926 20364 14960 20398
rect 14926 20296 14960 20326
rect 14926 20228 14960 20254
rect 14926 20160 14960 20182
rect 14926 20092 14960 20110
rect 14926 20024 14960 20038
rect 14926 19956 14960 19966
rect 14926 19888 14960 19894
rect 14926 19820 14960 19822
rect 14926 19784 14960 19786
rect 14926 19712 14960 19718
rect 14926 19640 14960 19650
rect 14926 19568 14960 19582
rect 14926 19496 14960 19514
rect 14926 19424 14960 19446
rect 14926 19352 14960 19378
rect 14716 19280 14870 19300
rect 14716 19276 14830 19280
rect 14750 19242 14830 19276
rect 14864 19242 14870 19280
rect 14716 19208 14870 19242
rect 14750 19174 14830 19208
rect 14864 19174 14870 19208
rect 14716 19170 14870 19174
rect 14926 19280 14960 19310
rect 14926 19208 14960 19242
rect 14716 19140 14750 19170
rect 14830 19156 14864 19170
rect 14926 19156 14960 19174
rect 15022 20432 15056 20450
rect 15022 20364 15056 20398
rect 15022 20296 15056 20326
rect 15022 20228 15056 20254
rect 15022 20160 15056 20182
rect 15022 20092 15056 20110
rect 15022 20024 15056 20038
rect 15022 19956 15056 19966
rect 15022 19888 15056 19894
rect 15022 19820 15056 19822
rect 15022 19784 15056 19786
rect 15022 19712 15056 19718
rect 15022 19640 15056 19650
rect 15022 19568 15056 19582
rect 15022 19496 15056 19514
rect 15022 19424 15056 19446
rect 15022 19352 15056 19378
rect 15022 19280 15056 19310
rect 15022 19208 15056 19242
rect 15022 19156 15056 19174
rect 15118 20432 15152 20450
rect 15118 20364 15152 20398
rect 15118 20296 15152 20326
rect 15118 20228 15152 20254
rect 15118 20160 15152 20182
rect 15118 20092 15152 20110
rect 15118 20024 15152 20038
rect 15118 19956 15152 19966
rect 15118 19888 15152 19894
rect 15118 19820 15152 19822
rect 15118 19784 15152 19786
rect 15118 19712 15152 19718
rect 15118 19640 15152 19650
rect 15118 19568 15152 19582
rect 15118 19496 15152 19514
rect 15118 19424 15152 19446
rect 15118 19352 15152 19378
rect 15118 19280 15152 19310
rect 15118 19208 15152 19242
rect 15118 19156 15152 19174
rect 15214 20432 15248 20450
rect 15214 20364 15248 20398
rect 15214 20296 15248 20326
rect 15214 20228 15248 20254
rect 15214 20160 15248 20182
rect 15214 20092 15248 20110
rect 15214 20024 15248 20038
rect 15214 19956 15248 19966
rect 15214 19888 15248 19894
rect 15214 19820 15248 19822
rect 15214 19784 15248 19786
rect 15214 19712 15248 19718
rect 15214 19640 15248 19650
rect 15214 19568 15248 19582
rect 15214 19496 15248 19514
rect 15214 19424 15248 19446
rect 15214 19352 15248 19378
rect 15214 19280 15248 19310
rect 15214 19208 15248 19242
rect 15214 19156 15248 19174
rect 15310 20432 15344 20450
rect 15310 20364 15344 20398
rect 15310 20296 15344 20326
rect 15310 20228 15344 20254
rect 15310 20160 15344 20182
rect 15310 20092 15344 20110
rect 15310 20024 15344 20038
rect 15310 19956 15344 19966
rect 15310 19888 15344 19894
rect 15310 19820 15344 19822
rect 15310 19784 15344 19786
rect 15310 19712 15344 19718
rect 15310 19640 15344 19650
rect 15310 19568 15344 19582
rect 15310 19496 15344 19514
rect 15310 19424 15344 19446
rect 15310 19352 15344 19378
rect 15310 19280 15344 19310
rect 15310 19208 15344 19242
rect 15310 19156 15344 19174
rect 15406 20432 15440 20450
rect 15406 20364 15440 20398
rect 15406 20296 15440 20326
rect 15406 20228 15440 20254
rect 15406 20160 15440 20182
rect 15406 20092 15440 20110
rect 15406 20024 15440 20038
rect 15406 19956 15440 19966
rect 15406 19888 15440 19894
rect 15406 19820 15440 19822
rect 15406 19784 15440 19786
rect 15406 19712 15440 19718
rect 15406 19640 15440 19650
rect 15406 19568 15440 19582
rect 15406 19496 15440 19514
rect 15406 19424 15440 19446
rect 15406 19352 15440 19378
rect 15406 19280 15440 19310
rect 15406 19208 15440 19242
rect 15406 19156 15440 19174
rect 15502 20432 15536 20450
rect 15502 20364 15536 20398
rect 15502 20296 15536 20326
rect 15502 20228 15536 20254
rect 15502 20160 15536 20182
rect 15502 20092 15536 20110
rect 15502 20024 15536 20038
rect 15502 19956 15536 19966
rect 15502 19888 15536 19894
rect 15502 19820 15536 19822
rect 15502 19784 15536 19786
rect 15502 19712 15536 19718
rect 15502 19640 15536 19650
rect 15502 19568 15536 19582
rect 15502 19496 15536 19514
rect 15502 19424 15536 19446
rect 15502 19352 15536 19378
rect 15502 19280 15536 19310
rect 15502 19208 15536 19242
rect 15502 19156 15536 19174
rect 15616 20432 15650 20466
rect 15616 20364 15650 20398
rect 15616 20296 15650 20330
rect 15616 20228 15650 20262
rect 15616 20160 15650 20194
rect 16656 20611 16690 20645
rect 16656 20543 16690 20577
rect 16656 20475 16690 20509
rect 16656 20407 16690 20441
rect 16656 20339 16690 20373
rect 16656 20271 16690 20305
rect 16656 20203 16690 20237
rect 16656 20135 16690 20169
rect 15616 20092 15650 20126
rect 15616 20024 15650 20058
rect 15616 19956 15650 19990
rect 15616 19888 15650 19922
rect 15616 19820 15650 19854
rect 15616 19752 15650 19786
rect 15616 19684 15650 19718
rect 15616 19616 15650 19650
rect 15616 19548 15650 19582
rect 15616 19480 15650 19514
rect 15616 19412 15650 19446
rect 15616 19344 15650 19378
rect 15616 19276 15650 19310
rect 15616 19208 15650 19242
rect 15616 19140 15650 19174
rect 14716 19020 14750 19106
rect 14862 19088 14878 19122
rect 14912 19088 14928 19122
rect 15054 19088 15070 19122
rect 15104 19088 15120 19122
rect 15246 19088 15262 19122
rect 15296 19088 15312 19122
rect 15438 19088 15454 19122
rect 15488 19088 15504 19122
rect 15616 19020 15650 19106
rect 14716 18986 14826 19020
rect 14860 18986 14894 19020
rect 14928 18986 14962 19020
rect 14996 18986 15030 19020
rect 15064 18986 15098 19020
rect 15132 18986 15166 19020
rect 15200 18986 15234 19020
rect 15268 18986 15302 19020
rect 15336 18986 15370 19020
rect 15404 18986 15438 19020
rect 15472 18986 15506 19020
rect 15540 18986 15650 19020
rect 15876 20100 15998 20134
rect 16032 20100 16066 20134
rect 16100 20100 16134 20134
rect 16168 20100 16202 20134
rect 16236 20100 16270 20134
rect 16304 20100 16426 20134
rect 15876 20019 15910 20100
rect 16118 19998 16134 20032
rect 16168 19998 16184 20032
rect 16392 20019 16426 20100
rect 15876 19951 15910 19985
rect 15876 19883 15910 19917
rect 15876 19815 15910 19849
rect 15876 19747 15910 19781
rect 15876 19679 15910 19713
rect 15876 19611 15910 19645
rect 15876 19543 15910 19577
rect 15876 19475 15910 19509
rect 15876 19407 15910 19441
rect 15876 19339 15910 19373
rect 15876 19271 15910 19305
rect 15876 19203 15910 19237
rect 15876 19135 15910 19169
rect 15990 19937 16024 19964
rect 15990 19865 16024 19883
rect 15990 19793 16024 19815
rect 15990 19721 16024 19747
rect 15990 19649 16024 19679
rect 15990 19577 16024 19611
rect 15990 19509 16024 19543
rect 15990 19441 16024 19471
rect 15990 19373 16024 19399
rect 15990 19305 16024 19327
rect 15990 19237 16024 19255
rect 15990 19156 16024 19183
rect 16086 19937 16120 19964
rect 16086 19865 16120 19883
rect 16086 19793 16120 19815
rect 16086 19721 16120 19747
rect 16086 19649 16120 19679
rect 16086 19577 16120 19611
rect 16086 19509 16120 19543
rect 16086 19441 16120 19471
rect 16086 19373 16120 19399
rect 16086 19305 16120 19327
rect 16086 19237 16120 19255
rect 16086 19156 16120 19183
rect 16182 19937 16216 19964
rect 16182 19865 16216 19883
rect 16182 19793 16216 19815
rect 16182 19721 16216 19747
rect 16182 19649 16216 19679
rect 16182 19577 16216 19611
rect 16182 19509 16216 19543
rect 16182 19441 16216 19471
rect 16182 19373 16216 19399
rect 16182 19305 16216 19327
rect 16182 19237 16216 19255
rect 16182 19156 16216 19183
rect 16278 19937 16312 19964
rect 16278 19865 16312 19883
rect 16278 19793 16312 19815
rect 16278 19721 16312 19747
rect 16278 19649 16312 19679
rect 16278 19577 16312 19611
rect 16278 19509 16312 19543
rect 16278 19441 16312 19471
rect 16278 19373 16312 19399
rect 16278 19305 16312 19327
rect 16278 19237 16312 19255
rect 16278 19156 16312 19183
rect 16392 19951 16426 19985
rect 16392 19883 16426 19917
rect 16392 19815 16426 19849
rect 16392 19747 16426 19781
rect 16392 19679 16426 19713
rect 16392 19611 16426 19645
rect 16392 19543 16426 19577
rect 16392 19475 16426 19509
rect 16392 19407 16426 19441
rect 16392 19339 16426 19373
rect 16392 19271 16426 19305
rect 16392 19203 16426 19237
rect 16392 19135 16426 19169
rect 15876 19020 15910 19101
rect 16022 19088 16038 19122
rect 16072 19088 16088 19122
rect 16214 19088 16230 19122
rect 16264 19088 16280 19122
rect 16392 19020 16426 19101
rect 15876 18986 15998 19020
rect 16032 18986 16066 19020
rect 16100 18986 16134 19020
rect 16168 18986 16202 19020
rect 16236 18986 16270 19020
rect 16304 18986 16426 19020
rect 16656 20067 16690 20101
rect 16656 19999 16690 20033
rect 16656 19931 16690 19965
rect 16656 19863 16690 19897
rect 16656 19795 16690 19829
rect 16656 19727 16690 19761
rect 16656 19659 16690 19693
rect 16656 19591 16690 19625
rect 16656 19523 16690 19557
rect 16656 19455 16690 19489
rect 16656 19387 16690 19421
rect 16656 19319 16690 19353
rect 16952 20883 16986 20917
rect 16952 20815 16986 20849
rect 16952 20747 16986 20781
rect 16952 20679 16986 20713
rect 16952 20611 16986 20645
rect 16952 20543 16986 20577
rect 16952 20475 16986 20509
rect 16952 20407 16986 20441
rect 16952 20339 16986 20373
rect 16952 20271 16986 20305
rect 16952 20203 16986 20237
rect 16952 20135 16986 20169
rect 16952 20067 16986 20101
rect 16952 19999 16986 20033
rect 16952 19931 16986 19965
rect 16952 19863 16986 19897
rect 16952 19795 16986 19829
rect 16952 19727 16986 19761
rect 16952 19659 16986 19693
rect 16952 19591 16986 19625
rect 16952 19523 16986 19557
rect 16952 19455 16986 19489
rect 16952 19387 16986 19421
rect 16952 19319 16986 19353
rect 16656 19251 16690 19285
rect 16656 19183 16690 19217
rect 16656 19115 16690 19149
rect 16656 19047 16690 19081
rect 13182 18871 13216 18905
rect 13182 18803 13216 18837
rect 14410 18939 14444 18973
rect 14410 18871 14444 18905
rect 13182 18735 13216 18769
rect 13182 18667 13216 18701
rect 13182 18599 13216 18633
rect 14410 18803 14444 18837
rect 14410 18735 14444 18769
rect 16656 18979 16690 19013
rect 16656 18911 16690 18945
rect 16952 19251 16986 19285
rect 16952 19183 16986 19217
rect 16952 19115 16986 19149
rect 16952 19047 16986 19081
rect 16952 18979 16986 19013
rect 16952 18911 16986 18945
rect 16656 18790 16690 18877
rect 16952 18790 16986 18877
rect 16656 18756 16770 18790
rect 16804 18756 16838 18790
rect 16872 18756 16986 18790
rect 17020 19232 17230 21565
rect 17020 19198 17072 19232
rect 17106 19198 17144 19232
rect 17178 19198 17230 19232
rect 14410 18667 14444 18701
rect 14410 18599 14444 18633
rect 13182 18531 13216 18565
rect 13182 18463 13216 18497
rect 14410 18531 14444 18565
rect 14410 18463 14444 18497
rect 13182 18395 13216 18429
rect 13182 18327 13216 18361
rect 13182 18259 13216 18293
rect 13182 18191 13216 18225
rect 14410 18395 14444 18429
rect 14410 18327 14444 18361
rect 14410 18259 14444 18293
rect 14410 18191 14444 18225
rect 13182 18123 13216 18157
rect 13182 18055 13216 18089
rect 14410 18123 14444 18157
rect 14410 18055 14444 18089
rect 13182 17987 13216 18021
rect 13182 17919 13216 17953
rect 13182 17851 13216 17885
rect 13182 17783 13216 17817
rect 14410 17987 14444 18021
rect 14902 18634 15026 18668
rect 15060 18634 15094 18668
rect 15128 18634 15252 18668
rect 14902 18547 14936 18634
rect 15044 18532 15060 18566
rect 15094 18532 15110 18566
rect 15218 18547 15252 18634
rect 14902 18479 14936 18513
rect 14902 18411 14936 18445
rect 14902 18343 14936 18377
rect 14902 18275 14936 18309
rect 14902 18207 14936 18241
rect 14902 18139 14936 18173
rect 14902 18071 14936 18105
rect 14902 18003 14936 18037
rect 14410 17919 14444 17953
rect 14410 17851 14444 17885
rect 13182 17715 13216 17749
rect 13182 17647 13216 17681
rect 14410 17783 14444 17817
rect 14410 17715 14444 17749
rect 13182 17579 13216 17613
rect 13182 17511 13216 17545
rect 13182 17443 13216 17477
rect 14410 17647 14444 17681
rect 14410 17579 14444 17613
rect 14410 17511 14444 17545
rect 14410 17443 14444 17477
rect 13182 17375 13216 17409
rect 13182 17307 13216 17341
rect 14410 17375 14444 17409
rect 14410 17307 14444 17341
rect 13182 17239 13216 17273
rect 13182 17171 13216 17205
rect 13182 17103 13216 17137
rect 13182 17035 13216 17069
rect 14410 17239 14444 17273
rect 14410 17171 14444 17205
rect 14410 17103 14444 17137
rect 14410 17035 14444 17069
rect 13182 16967 13216 17001
rect 13182 16899 13216 16933
rect 14410 16967 14444 17001
rect 14410 16899 14444 16933
rect 13182 16794 13216 16865
rect 14410 16794 14444 16865
rect 13182 16760 13286 16794
rect 13320 16760 13354 16794
rect 13388 16760 13422 16794
rect 13456 16760 13490 16794
rect 13524 16760 13558 16794
rect 13592 16760 13626 16794
rect 13660 16760 13694 16794
rect 13728 16760 13762 16794
rect 13796 16760 13830 16794
rect 13864 16760 13898 16794
rect 13932 16760 13966 16794
rect 14000 16760 14034 16794
rect 14068 16760 14102 16794
rect 14136 16760 14170 16794
rect 14204 16760 14238 16794
rect 14272 16760 14306 16794
rect 14340 16760 14444 16794
rect 14512 17950 14626 17984
rect 14660 17950 14694 17984
rect 14728 17950 14842 17984
rect 14512 17865 14546 17950
rect 14808 17865 14842 17950
rect 14512 17797 14546 17831
rect 14512 17729 14546 17763
rect 14512 17661 14546 17695
rect 14512 17593 14546 17627
rect 14512 17525 14546 17559
rect 14512 17457 14546 17491
rect 14512 17389 14546 17423
rect 14808 17797 14842 17831
rect 14808 17729 14842 17763
rect 14808 17661 14842 17695
rect 14808 17593 14842 17627
rect 14808 17525 14842 17559
rect 14808 17457 14842 17491
rect 14512 17321 14546 17355
rect 14808 17389 14842 17423
rect 14512 17253 14546 17287
rect 14512 17185 14546 17219
rect 14512 17117 14546 17151
rect 14512 17049 14546 17083
rect 14512 16981 14546 17015
rect 14512 16913 14546 16947
rect 14808 17321 14842 17355
rect 14808 17253 14842 17287
rect 14808 17185 14842 17219
rect 14808 17117 14842 17151
rect 14808 17049 14842 17083
rect 14808 16981 14842 17015
rect 14808 16913 14842 16947
rect 14512 16794 14546 16879
rect 14808 16794 14842 16879
rect 14512 16760 14626 16794
rect 14660 16760 14694 16794
rect 14728 16760 14842 16794
rect 14902 17935 14936 17969
rect 14902 17867 14936 17901
rect 14902 17799 14936 17833
rect 14902 17731 14936 17765
rect 14902 17663 14936 17697
rect 14902 17595 14936 17629
rect 14902 17527 14936 17561
rect 14902 17459 14936 17493
rect 14902 17391 14936 17425
rect 14902 17323 14936 17357
rect 14902 17255 14936 17289
rect 14902 17187 14936 17221
rect 14902 17119 14936 17153
rect 14902 17051 14936 17085
rect 14902 16983 14936 17017
rect 14902 16915 14936 16949
rect 15016 18479 15050 18498
rect 15016 18411 15050 18417
rect 15016 18343 15050 18345
rect 15016 18307 15050 18309
rect 15016 18235 15050 18241
rect 15016 18163 15050 18173
rect 15016 18091 15050 18105
rect 15016 18019 15050 18037
rect 15016 17947 15050 17969
rect 15016 17875 15050 17901
rect 15016 17803 15050 17833
rect 15016 17731 15050 17765
rect 15016 17663 15050 17697
rect 15016 17595 15050 17625
rect 15016 17527 15050 17553
rect 15016 17459 15050 17481
rect 15016 17391 15050 17409
rect 15016 17323 15050 17337
rect 15016 17255 15050 17265
rect 15016 17187 15050 17193
rect 15016 17119 15050 17121
rect 15016 17083 15050 17085
rect 15016 17011 15050 17017
rect 15016 16930 15050 16949
rect 15104 18479 15138 18498
rect 15104 18411 15138 18417
rect 15104 18343 15138 18345
rect 15104 18307 15138 18309
rect 15104 18235 15138 18241
rect 15104 18163 15138 18173
rect 15104 18091 15138 18105
rect 15104 18019 15138 18037
rect 15104 17947 15138 17969
rect 15104 17875 15138 17901
rect 15104 17803 15138 17833
rect 15104 17731 15138 17765
rect 15104 17663 15138 17697
rect 15104 17595 15138 17625
rect 15104 17527 15138 17553
rect 15104 17459 15138 17481
rect 15104 17391 15138 17409
rect 15104 17323 15138 17337
rect 15104 17255 15138 17265
rect 15104 17187 15138 17193
rect 15104 17119 15138 17121
rect 15104 17083 15138 17085
rect 15104 17011 15138 17017
rect 15104 16930 15138 16949
rect 15218 18479 15252 18513
rect 15218 18411 15252 18445
rect 15218 18343 15252 18377
rect 15312 18634 15436 18668
rect 15470 18634 15504 18668
rect 15538 18634 15662 18668
rect 15312 18547 15346 18634
rect 15454 18532 15470 18566
rect 15504 18532 15520 18566
rect 15628 18547 15662 18634
rect 15312 18479 15346 18513
rect 15312 18411 15346 18445
rect 15312 18343 15346 18377
rect 15218 18275 15252 18309
rect 15218 18207 15252 18241
rect 15218 18139 15252 18173
rect 15218 18071 15252 18105
rect 15308 18309 15312 18329
rect 15426 18479 15460 18498
rect 15426 18411 15460 18417
rect 15426 18343 15460 18345
rect 15346 18309 15426 18329
rect 15308 18307 15460 18309
rect 15308 18275 15426 18307
rect 15308 18241 15312 18275
rect 15346 18241 15426 18275
rect 15308 18235 15460 18241
rect 15308 18207 15426 18235
rect 15308 18173 15312 18207
rect 15346 18173 15426 18207
rect 15308 18163 15460 18173
rect 15308 18139 15426 18163
rect 15308 18105 15312 18139
rect 15346 18105 15426 18139
rect 15308 18091 15460 18105
rect 15308 18077 15426 18091
rect 15218 18003 15252 18037
rect 15218 17935 15252 17969
rect 15218 17867 15252 17901
rect 15218 17799 15252 17833
rect 15218 17731 15252 17765
rect 15218 17663 15252 17697
rect 15218 17595 15252 17629
rect 15218 17527 15252 17561
rect 15218 17459 15252 17493
rect 15218 17391 15252 17425
rect 15218 17323 15252 17357
rect 15218 17255 15252 17289
rect 15218 17187 15252 17221
rect 15218 17119 15252 17153
rect 15218 17051 15252 17085
rect 15218 16983 15252 17017
rect 15218 16915 15252 16949
rect 14902 16794 14936 16881
rect 15044 16862 15060 16896
rect 15094 16862 15110 16896
rect 15218 16794 15252 16881
rect 14902 16760 15026 16794
rect 15060 16760 15094 16794
rect 15128 16760 15252 16794
rect 15312 18071 15346 18077
rect 15312 18003 15346 18037
rect 15312 17935 15346 17969
rect 15312 17867 15346 17901
rect 15312 17799 15346 17833
rect 15312 17731 15346 17765
rect 15312 17663 15346 17697
rect 15312 17595 15346 17629
rect 15312 17527 15346 17561
rect 15312 17459 15346 17493
rect 15312 17391 15346 17425
rect 15312 17323 15346 17357
rect 15312 17255 15346 17289
rect 15312 17187 15346 17221
rect 15312 17119 15346 17153
rect 15312 17051 15346 17085
rect 15312 16983 15346 17017
rect 15312 16915 15346 16949
rect 15426 18019 15460 18037
rect 15426 17947 15460 17969
rect 15426 17875 15460 17901
rect 15426 17803 15460 17833
rect 15426 17731 15460 17765
rect 15426 17663 15460 17697
rect 15426 17595 15460 17625
rect 15426 17527 15460 17553
rect 15426 17459 15460 17481
rect 15426 17391 15460 17409
rect 15426 17323 15460 17337
rect 15426 17255 15460 17265
rect 15426 17187 15460 17193
rect 15426 17119 15460 17121
rect 15426 17083 15460 17085
rect 15426 17011 15460 17017
rect 15426 16930 15460 16949
rect 15514 18479 15548 18498
rect 15514 18411 15548 18417
rect 15514 18343 15548 18345
rect 15514 18307 15548 18309
rect 15514 18235 15548 18241
rect 15514 18163 15548 18173
rect 15514 18091 15548 18105
rect 15514 18019 15548 18037
rect 15514 17947 15548 17969
rect 15514 17875 15548 17901
rect 15514 17803 15548 17833
rect 15514 17731 15548 17765
rect 15514 17663 15548 17697
rect 15514 17595 15548 17625
rect 15514 17527 15548 17553
rect 15514 17459 15548 17481
rect 15514 17391 15548 17409
rect 15514 17323 15548 17337
rect 15514 17255 15548 17265
rect 15514 17187 15548 17193
rect 15514 17119 15548 17121
rect 15514 17083 15548 17085
rect 15514 17011 15548 17017
rect 15514 16930 15548 16949
rect 15628 18479 15662 18513
rect 15628 18411 15662 18445
rect 15628 18343 15662 18377
rect 15628 18275 15662 18309
rect 15628 18207 15662 18241
rect 15628 18139 15662 18173
rect 15628 18071 15662 18105
rect 15628 18003 15662 18037
rect 16124 18651 16238 18685
rect 16272 18651 16306 18685
rect 16340 18651 16454 18685
rect 16124 18556 16158 18651
rect 16420 18556 16454 18651
rect 16124 18488 16158 18522
rect 16124 18420 16158 18454
rect 16124 18352 16158 18386
rect 16124 18284 16158 18318
rect 16124 18216 16158 18250
rect 16124 18148 16158 18182
rect 16420 18488 16454 18522
rect 16750 18460 16910 18756
rect 16420 18420 16454 18454
rect 16420 18352 16454 18386
rect 16420 18284 16454 18318
rect 16420 18216 16454 18250
rect 16420 18148 16454 18182
rect 16686 18426 16782 18460
rect 16816 18426 16850 18460
rect 16884 18426 16980 18460
rect 16686 18364 16720 18426
rect 16946 18364 16980 18426
rect 16686 18296 16720 18330
rect 16784 18330 16882 18346
rect 16784 18296 16816 18330
rect 16850 18296 16882 18330
rect 16784 18280 16882 18296
rect 16946 18296 16980 18330
rect 16686 18200 16720 18262
rect 16946 18200 16980 18262
rect 16686 18166 16782 18200
rect 16816 18166 16850 18200
rect 16884 18166 16980 18200
rect 16124 18080 16158 18114
rect 16124 18012 16158 18046
rect 15628 17935 15662 17969
rect 15628 17867 15662 17901
rect 15628 17799 15662 17833
rect 15628 17731 15662 17765
rect 15628 17663 15662 17697
rect 15628 17595 15662 17629
rect 15628 17527 15662 17561
rect 15628 17459 15662 17493
rect 15628 17391 15662 17425
rect 15628 17323 15662 17357
rect 15628 17255 15662 17289
rect 15628 17187 15662 17221
rect 15628 17119 15662 17153
rect 15628 17051 15662 17085
rect 15628 16983 15662 17017
rect 15628 16915 15662 16949
rect 15312 16794 15346 16881
rect 15454 16862 15470 16896
rect 15504 16862 15520 16896
rect 15628 16794 15662 16881
rect 15312 16760 15436 16794
rect 15470 16760 15504 16794
rect 15538 16760 15662 16794
rect 15732 17950 15846 17984
rect 15880 17950 15914 17984
rect 15948 17950 16062 17984
rect 15732 17865 15766 17950
rect 16028 17865 16062 17950
rect 15732 17797 15766 17831
rect 15732 17729 15766 17763
rect 15732 17661 15766 17695
rect 15732 17593 15766 17627
rect 15732 17525 15766 17559
rect 15732 17457 15766 17491
rect 15732 17389 15766 17423
rect 16028 17797 16062 17831
rect 16028 17729 16062 17763
rect 16028 17661 16062 17695
rect 16028 17593 16062 17627
rect 16028 17525 16062 17559
rect 16028 17457 16062 17491
rect 15732 17321 15766 17355
rect 16028 17389 16062 17423
rect 15732 17253 15766 17287
rect 15732 17185 15766 17219
rect 15732 17117 15766 17151
rect 15732 17049 15766 17083
rect 15732 16981 15766 17015
rect 15732 16913 15766 16947
rect 16028 17321 16062 17355
rect 16028 17253 16062 17287
rect 16028 17185 16062 17219
rect 16028 17117 16062 17151
rect 16028 17049 16062 17083
rect 16028 16981 16062 17015
rect 16028 16913 16062 16947
rect 15732 16794 15766 16879
rect 16028 16794 16062 16879
rect 15732 16760 15846 16794
rect 15880 16760 15914 16794
rect 15948 16760 16062 16794
rect 16124 17944 16158 17978
rect 16124 17876 16158 17910
rect 16124 17808 16158 17842
rect 16124 17740 16158 17774
rect 16124 17672 16158 17706
rect 16124 17604 16158 17638
rect 16124 17536 16158 17570
rect 16124 17468 16158 17502
rect 16124 17400 16158 17434
rect 16124 17332 16158 17366
rect 16420 18080 16454 18114
rect 16420 18012 16454 18046
rect 16420 17944 16454 17978
rect 16420 17876 16454 17910
rect 16420 17808 16454 17842
rect 16420 17740 16454 17774
rect 16420 17672 16454 17706
rect 16420 17604 16454 17638
rect 16420 17536 16454 17570
rect 16420 17468 16454 17502
rect 16420 17400 16454 17434
rect 16420 17332 16454 17366
rect 16124 17264 16158 17298
rect 16124 17196 16158 17230
rect 16124 17128 16158 17162
rect 16124 17060 16158 17094
rect 16124 16992 16158 17026
rect 16124 16924 16158 16958
rect 16420 17264 16454 17298
rect 16420 17196 16454 17230
rect 16420 17128 16454 17162
rect 16420 17060 16454 17094
rect 16420 16992 16454 17026
rect 16420 16924 16454 16958
rect 16124 16795 16158 16890
rect 16420 16795 16454 16890
rect 16124 16761 16238 16795
rect 16272 16761 16306 16795
rect 16340 16761 16454 16795
rect 17020 17280 17230 19198
rect 17266 21466 17380 21500
rect 17414 21466 17448 21500
rect 17482 21466 17596 21500
rect 17266 21393 17300 21466
rect 17562 21393 17596 21466
rect 17266 21325 17300 21359
rect 17266 21257 17300 21291
rect 17266 21189 17300 21223
rect 17266 21121 17300 21155
rect 17266 21053 17300 21087
rect 17266 20985 17300 21019
rect 17266 20917 17300 20951
rect 17562 21325 17596 21359
rect 17562 21257 17596 21291
rect 17562 21189 17596 21223
rect 17562 21121 17596 21155
rect 17562 21053 17596 21087
rect 17562 20985 17596 21019
rect 17266 20849 17300 20883
rect 17266 20781 17300 20815
rect 17266 20713 17300 20747
rect 17266 20645 17300 20679
rect 17266 20577 17300 20611
rect 17266 20509 17300 20543
rect 17266 20441 17300 20475
rect 17266 20373 17300 20407
rect 17266 20305 17300 20339
rect 17266 20237 17300 20271
rect 17266 20169 17300 20203
rect 17266 20101 17300 20135
rect 17266 20033 17300 20067
rect 17266 19965 17300 19999
rect 17266 19897 17300 19931
rect 17266 19829 17300 19863
rect 17266 19761 17300 19795
rect 17266 19693 17300 19727
rect 17266 19625 17300 19659
rect 17266 19557 17300 19591
rect 17266 19489 17300 19523
rect 17266 19421 17300 19455
rect 17266 19353 17300 19387
rect 17266 19285 17300 19319
rect 17266 19217 17300 19251
rect 17266 19149 17300 19183
rect 17266 19081 17300 19115
rect 17266 19013 17300 19047
rect 17266 18945 17300 18979
rect 17266 18877 17300 18911
rect 17266 18809 17300 18843
rect 17266 18741 17300 18775
rect 17266 18673 17300 18707
rect 17266 18605 17300 18639
rect 17266 18537 17300 18571
rect 17266 18469 17300 18503
rect 17266 18401 17300 18435
rect 17266 18333 17300 18367
rect 17266 18265 17300 18299
rect 17266 18197 17300 18231
rect 17266 18129 17300 18163
rect 17266 18061 17300 18095
rect 17266 17993 17300 18027
rect 17266 17925 17300 17959
rect 17562 20917 17596 20951
rect 17562 20849 17596 20883
rect 17562 20781 17596 20815
rect 17562 20713 17596 20747
rect 17562 20645 17596 20679
rect 17562 20577 17596 20611
rect 17562 20509 17596 20543
rect 17562 20441 17596 20475
rect 17562 20373 17596 20407
rect 17562 20305 17596 20339
rect 17562 20237 17596 20271
rect 17562 20169 17596 20203
rect 17562 20101 17596 20135
rect 17562 20033 17596 20067
rect 17562 19965 17596 19999
rect 17562 19897 17596 19931
rect 17562 19829 17596 19863
rect 17562 19761 17596 19795
rect 17562 19693 17596 19727
rect 17562 19625 17596 19659
rect 17562 19557 17596 19591
rect 17562 19489 17596 19523
rect 17562 19421 17596 19455
rect 17562 19353 17596 19387
rect 17562 19285 17596 19319
rect 17562 19217 17596 19251
rect 17562 19149 17596 19183
rect 17562 19081 17596 19115
rect 17562 19013 17596 19047
rect 17562 18945 17596 18979
rect 17562 18877 17596 18911
rect 17562 18809 17596 18843
rect 17562 18741 17596 18775
rect 17562 18673 17596 18707
rect 17562 18605 17596 18639
rect 17562 18537 17596 18571
rect 17562 18469 17596 18503
rect 17562 18401 17596 18435
rect 17562 18333 17596 18367
rect 17562 18265 17596 18299
rect 17562 18197 17596 18231
rect 17562 18129 17596 18163
rect 17562 18061 17596 18095
rect 17562 17993 17596 18027
rect 17266 17857 17300 17891
rect 17266 17789 17300 17823
rect 17266 17721 17300 17755
rect 17266 17653 17300 17687
rect 17266 17585 17300 17619
rect 17266 17517 17300 17551
rect 17562 17925 17596 17959
rect 17562 17857 17596 17891
rect 17562 17789 17596 17823
rect 17562 17721 17596 17755
rect 17562 17653 17596 17687
rect 17562 17585 17596 17619
rect 17562 17517 17596 17551
rect 17266 17410 17300 17483
rect 17562 17410 17596 17483
rect 17266 17376 17380 17410
rect 17414 17376 17448 17410
rect 17482 17376 17596 17410
rect 17020 16460 17240 17280
rect 13306 16432 17240 16460
rect 13306 16326 13338 16432
rect 13444 16401 17240 16432
rect 13444 16367 14623 16401
rect 14657 16367 14695 16401
rect 14729 16367 15838 16401
rect 15872 16367 15910 16401
rect 15944 16367 17240 16401
rect 13444 16326 17240 16367
rect 13306 16308 17240 16326
rect 16941 16245 17240 16308
rect 16941 16140 17561 16245
rect 16940 16126 17561 16140
rect 14308 16044 14432 16078
rect 14466 16044 14500 16078
rect 14534 16044 14568 16078
rect 14602 16044 14636 16078
rect 14670 16044 14704 16078
rect 14738 16044 14772 16078
rect 14806 16044 14840 16078
rect 14874 16044 14908 16078
rect 14942 16044 14976 16078
rect 15010 16044 15044 16078
rect 15078 16044 15112 16078
rect 15146 16044 15180 16078
rect 15214 16044 15338 16078
rect 14308 15975 14342 16044
rect 14550 15942 14566 15976
rect 14600 15942 14616 15976
rect 14742 15942 14758 15976
rect 14792 15942 14808 15976
rect 14934 15942 14950 15976
rect 14984 15942 15000 15976
rect 15126 15942 15142 15976
rect 15176 15942 15192 15976
rect 15304 15975 15338 16044
rect 14308 15907 14342 15941
rect 14308 15839 14342 15873
rect 14308 15771 14342 15805
rect 14308 15703 14342 15737
rect 13458 15604 13582 15638
rect 13616 15604 13650 15638
rect 13684 15604 13808 15638
rect 13458 15517 13492 15604
rect 13600 15502 13616 15536
rect 13650 15502 13666 15536
rect 13774 15517 13808 15604
rect 13458 15449 13492 15483
rect 13458 15381 13492 15415
rect 13458 15313 13492 15347
rect 13458 15245 13492 15279
rect 13458 15177 13492 15211
rect 13458 15109 13492 15143
rect 13458 15041 13492 15075
rect 13458 14973 13492 15007
rect 13458 14905 13492 14939
rect 13458 14837 13492 14871
rect 13458 14769 13492 14803
rect 13458 14701 13492 14735
rect 13458 14633 13492 14667
rect 13458 14565 13492 14599
rect 13458 14497 13492 14531
rect 13458 14429 13492 14463
rect 13458 14361 13492 14395
rect 13458 14293 13492 14327
rect 13458 14225 13492 14259
rect 13458 14157 13492 14191
rect 13458 14089 13492 14123
rect 13458 14021 13492 14055
rect 13458 13953 13492 13987
rect 13458 13885 13492 13919
rect 13572 15449 13606 15468
rect 13660 15463 13694 15468
rect 13774 15463 13808 15483
rect 13572 15381 13606 15387
rect 13659 15449 13808 15463
rect 13659 15387 13660 15449
rect 13694 15415 13774 15449
rect 13694 15387 13808 15415
rect 13659 15381 13808 15387
rect 13659 15327 13660 15381
rect 13694 15347 13774 15381
rect 13572 15313 13606 15315
rect 13572 15277 13606 15279
rect 13572 15205 13606 15211
rect 13572 15133 13606 15143
rect 13572 15061 13606 15075
rect 13572 14989 13606 15007
rect 13572 14917 13606 14939
rect 13572 14845 13606 14871
rect 13572 14773 13606 14803
rect 13572 14701 13606 14735
rect 13572 14633 13606 14667
rect 13572 14565 13606 14595
rect 13572 14497 13606 14523
rect 13572 14429 13606 14451
rect 13572 14361 13606 14379
rect 13572 14293 13606 14307
rect 13572 14225 13606 14235
rect 13572 14157 13606 14163
rect 13572 14089 13606 14091
rect 13572 14053 13606 14055
rect 13572 13981 13606 13987
rect 13572 13900 13606 13919
rect 13694 15327 13808 15347
rect 13660 15313 13694 15315
rect 13660 15277 13694 15279
rect 13660 15205 13694 15211
rect 13660 15133 13694 15143
rect 13660 15061 13694 15075
rect 13660 14989 13694 15007
rect 13660 14917 13694 14939
rect 13660 14845 13694 14871
rect 13660 14773 13694 14803
rect 13660 14701 13694 14735
rect 13660 14633 13694 14667
rect 13660 14565 13694 14595
rect 13660 14497 13694 14523
rect 13660 14429 13694 14451
rect 13660 14361 13694 14379
rect 13660 14293 13694 14307
rect 13660 14225 13694 14235
rect 13660 14157 13694 14163
rect 13660 14089 13694 14091
rect 13660 14053 13694 14055
rect 13660 13981 13694 13987
rect 13660 13900 13694 13919
rect 13774 15313 13808 15327
rect 13774 15245 13808 15279
rect 13774 15177 13808 15211
rect 13774 15109 13808 15143
rect 13774 15041 13808 15075
rect 13774 14973 13808 15007
rect 13774 14905 13808 14939
rect 13774 14837 13808 14871
rect 13774 14769 13808 14803
rect 13774 14701 13808 14735
rect 13774 14633 13808 14667
rect 13774 14565 13808 14599
rect 13774 14497 13808 14531
rect 13774 14429 13808 14463
rect 13774 14361 13808 14395
rect 13774 14293 13808 14327
rect 13774 14225 13808 14259
rect 13774 14157 13808 14191
rect 13774 14089 13808 14123
rect 13774 14021 13808 14055
rect 13774 13953 13808 13987
rect 13774 13885 13808 13919
rect 13458 13764 13492 13851
rect 13600 13832 13616 13866
rect 13650 13832 13666 13866
rect 13774 13764 13808 13851
rect 13458 13730 13582 13764
rect 13616 13730 13650 13764
rect 13684 13730 13808 13764
rect 14308 15635 14342 15669
rect 14308 15567 14342 15601
rect 14308 15499 14342 15533
rect 14308 15431 14342 15465
rect 14308 15363 14342 15397
rect 14308 15295 14342 15329
rect 14308 15227 14342 15261
rect 14308 15159 14342 15193
rect 14308 15091 14342 15125
rect 14308 15023 14342 15057
rect 14308 14955 14342 14989
rect 14308 14887 14342 14921
rect 14308 14819 14342 14853
rect 14308 14751 14342 14785
rect 14308 14683 14342 14717
rect 14308 14615 14342 14649
rect 14308 14547 14342 14581
rect 14308 14479 14342 14513
rect 14308 14411 14342 14445
rect 14308 14343 14342 14377
rect 14308 14275 14342 14309
rect 14308 14207 14342 14241
rect 14308 14139 14342 14173
rect 14308 14071 14342 14105
rect 14308 14003 14342 14037
rect 14308 13935 14342 13969
rect 14308 13867 14342 13901
rect 14422 15873 14456 15908
rect 14422 15805 14456 15823
rect 14422 15737 14456 15751
rect 14422 15669 14456 15679
rect 14422 15601 14456 15607
rect 14422 15533 14456 15535
rect 14422 15497 14456 15499
rect 14422 15425 14456 15431
rect 14422 15353 14456 15363
rect 14422 15281 14456 15295
rect 14422 15209 14456 15227
rect 14422 15137 14456 15159
rect 14422 15065 14456 15091
rect 14422 14993 14456 15023
rect 14422 14921 14456 14955
rect 14422 14853 14456 14887
rect 14422 14785 14456 14815
rect 14422 14717 14456 14743
rect 14422 14649 14456 14671
rect 14422 14581 14456 14599
rect 14422 14513 14456 14527
rect 14422 14445 14456 14455
rect 14422 14377 14456 14383
rect 14422 14309 14456 14311
rect 14422 14273 14456 14275
rect 14422 14201 14456 14207
rect 14422 14129 14456 14139
rect 14422 14057 14456 14071
rect 14422 13985 14456 14003
rect 14422 13900 14456 13935
rect 14518 15873 14552 15908
rect 14518 15805 14552 15823
rect 14518 15737 14552 15751
rect 14518 15669 14552 15679
rect 14518 15601 14552 15607
rect 14518 15533 14552 15535
rect 14518 15497 14552 15499
rect 14518 15425 14552 15431
rect 14518 15353 14552 15363
rect 14518 15281 14552 15295
rect 14518 15209 14552 15227
rect 14518 15137 14552 15159
rect 14518 15065 14552 15091
rect 14518 14993 14552 15023
rect 14518 14921 14552 14955
rect 14518 14853 14552 14887
rect 14518 14785 14552 14815
rect 14518 14717 14552 14743
rect 14518 14649 14552 14671
rect 14518 14581 14552 14599
rect 14518 14513 14552 14527
rect 14518 14445 14552 14455
rect 14518 14377 14552 14383
rect 14518 14309 14552 14311
rect 14518 14273 14552 14275
rect 14518 14201 14552 14207
rect 14518 14129 14552 14139
rect 14518 14057 14552 14071
rect 14518 13985 14552 14003
rect 14518 13900 14552 13935
rect 14614 15873 14648 15908
rect 14614 15805 14648 15823
rect 14614 15737 14648 15751
rect 14614 15669 14648 15679
rect 14614 15601 14648 15607
rect 14614 15533 14648 15535
rect 14614 15497 14648 15499
rect 14614 15425 14648 15431
rect 14614 15353 14648 15363
rect 14614 15281 14648 15295
rect 14614 15209 14648 15227
rect 14614 15137 14648 15159
rect 14614 15065 14648 15091
rect 14614 14993 14648 15023
rect 14614 14921 14648 14955
rect 14614 14853 14648 14887
rect 14614 14785 14648 14815
rect 14614 14717 14648 14743
rect 14614 14649 14648 14671
rect 14614 14581 14648 14599
rect 14614 14513 14648 14527
rect 14614 14445 14648 14455
rect 14614 14377 14648 14383
rect 14614 14309 14648 14311
rect 14614 14273 14648 14275
rect 14614 14201 14648 14207
rect 14614 14129 14648 14139
rect 14614 14057 14648 14071
rect 14614 13985 14648 14003
rect 14614 13900 14648 13935
rect 14710 15873 14744 15908
rect 14710 15805 14744 15823
rect 14710 15737 14744 15751
rect 14710 15669 14744 15679
rect 14710 15601 14744 15607
rect 14710 15533 14744 15535
rect 14710 15497 14744 15499
rect 14710 15425 14744 15431
rect 14710 15353 14744 15363
rect 14710 15281 14744 15295
rect 14710 15209 14744 15227
rect 14710 15137 14744 15159
rect 14710 15065 14744 15091
rect 14710 14993 14744 15023
rect 14710 14921 14744 14955
rect 14710 14853 14744 14887
rect 14710 14785 14744 14815
rect 14710 14717 14744 14743
rect 14710 14649 14744 14671
rect 14710 14581 14744 14599
rect 14710 14513 14744 14527
rect 14710 14445 14744 14455
rect 14710 14377 14744 14383
rect 14710 14309 14744 14311
rect 14710 14273 14744 14275
rect 14710 14201 14744 14207
rect 14710 14129 14744 14139
rect 14710 14057 14744 14071
rect 14710 13985 14744 14003
rect 14710 13900 14744 13935
rect 14806 15873 14840 15908
rect 14806 15805 14840 15823
rect 14806 15737 14840 15751
rect 14806 15669 14840 15679
rect 14806 15601 14840 15607
rect 14806 15533 14840 15535
rect 14806 15497 14840 15499
rect 14806 15425 14840 15431
rect 14806 15353 14840 15363
rect 14806 15281 14840 15295
rect 14806 15209 14840 15227
rect 14806 15137 14840 15159
rect 14806 15065 14840 15091
rect 14806 14993 14840 15023
rect 14806 14921 14840 14955
rect 14806 14853 14840 14887
rect 14806 14785 14840 14815
rect 14806 14717 14840 14743
rect 14806 14649 14840 14671
rect 14806 14581 14840 14599
rect 14806 14513 14840 14527
rect 14806 14445 14840 14455
rect 14806 14377 14840 14383
rect 14806 14309 14840 14311
rect 14806 14273 14840 14275
rect 14806 14201 14840 14207
rect 14806 14129 14840 14139
rect 14806 14057 14840 14071
rect 14806 13985 14840 14003
rect 14806 13900 14840 13935
rect 14902 15873 14936 15908
rect 14902 15805 14936 15823
rect 14902 15737 14936 15751
rect 14902 15669 14936 15679
rect 14902 15601 14936 15607
rect 14902 15533 14936 15535
rect 14902 15497 14936 15499
rect 14902 15425 14936 15431
rect 14902 15353 14936 15363
rect 14902 15281 14936 15295
rect 14902 15209 14936 15227
rect 14902 15137 14936 15159
rect 14902 15065 14936 15091
rect 14902 14993 14936 15023
rect 14902 14921 14936 14955
rect 14902 14853 14936 14887
rect 14902 14785 14936 14815
rect 14902 14717 14936 14743
rect 14902 14649 14936 14671
rect 14902 14581 14936 14599
rect 14902 14513 14936 14527
rect 14902 14445 14936 14455
rect 14902 14377 14936 14383
rect 14902 14309 14936 14311
rect 14902 14273 14936 14275
rect 14902 14201 14936 14207
rect 14902 14129 14936 14139
rect 14902 14057 14936 14071
rect 14902 13985 14936 14003
rect 14902 13900 14936 13935
rect 14998 15873 15032 15908
rect 14998 15805 15032 15823
rect 14998 15737 15032 15751
rect 14998 15669 15032 15679
rect 14998 15601 15032 15607
rect 14998 15533 15032 15535
rect 14998 15497 15032 15499
rect 14998 15425 15032 15431
rect 14998 15353 15032 15363
rect 14998 15281 15032 15295
rect 14998 15209 15032 15227
rect 14998 15137 15032 15159
rect 14998 15065 15032 15091
rect 14998 14993 15032 15023
rect 14998 14921 15032 14955
rect 14998 14853 15032 14887
rect 14998 14785 15032 14815
rect 14998 14717 15032 14743
rect 14998 14649 15032 14671
rect 14998 14581 15032 14599
rect 14998 14513 15032 14527
rect 14998 14445 15032 14455
rect 14998 14377 15032 14383
rect 14998 14309 15032 14311
rect 14998 14273 15032 14275
rect 14998 14201 15032 14207
rect 14998 14129 15032 14139
rect 14998 14057 15032 14071
rect 14998 13985 15032 14003
rect 14998 13900 15032 13935
rect 15094 15873 15128 15908
rect 15094 15805 15128 15823
rect 15094 15737 15128 15751
rect 15094 15669 15128 15679
rect 15094 15601 15128 15607
rect 15094 15533 15128 15535
rect 15094 15497 15128 15499
rect 15094 15425 15128 15431
rect 15094 15353 15128 15363
rect 15094 15281 15128 15295
rect 15094 15209 15128 15227
rect 15094 15137 15128 15159
rect 15094 15065 15128 15091
rect 15094 14993 15128 15023
rect 15094 14921 15128 14955
rect 15094 14853 15128 14887
rect 15094 14785 15128 14815
rect 15094 14717 15128 14743
rect 15094 14649 15128 14671
rect 15094 14581 15128 14599
rect 15094 14513 15128 14527
rect 15094 14445 15128 14455
rect 15094 14377 15128 14383
rect 15094 14309 15128 14311
rect 15094 14273 15128 14275
rect 15094 14201 15128 14207
rect 15094 14129 15128 14139
rect 15094 14057 15128 14071
rect 15094 13985 15128 14003
rect 15094 13900 15128 13935
rect 15190 15873 15224 15908
rect 15190 15805 15224 15823
rect 15190 15737 15224 15751
rect 15190 15669 15224 15679
rect 15190 15601 15224 15607
rect 15190 15533 15224 15535
rect 15190 15497 15224 15499
rect 15190 15425 15224 15431
rect 15190 15353 15224 15363
rect 15190 15281 15224 15295
rect 15190 15209 15224 15227
rect 15190 15137 15224 15159
rect 15190 15065 15224 15091
rect 15190 14993 15224 15023
rect 15190 14921 15224 14955
rect 15190 14853 15224 14887
rect 15190 14785 15224 14815
rect 15190 14717 15224 14743
rect 15190 14649 15224 14671
rect 15190 14581 15224 14599
rect 15190 14513 15224 14527
rect 15190 14445 15224 14455
rect 15190 14377 15224 14383
rect 15190 14309 15224 14311
rect 15190 14273 15224 14275
rect 15190 14201 15224 14207
rect 15190 14129 15224 14139
rect 15190 14057 15224 14071
rect 15190 13985 15224 14003
rect 15190 13900 15224 13935
rect 15304 15907 15338 15941
rect 15304 15839 15338 15873
rect 15304 15771 15338 15805
rect 15304 15703 15338 15737
rect 15304 15635 15338 15669
rect 15304 15567 15338 15601
rect 15304 15499 15338 15533
rect 15304 15431 15338 15465
rect 15304 15363 15338 15397
rect 15304 15295 15338 15329
rect 15304 15227 15338 15261
rect 15304 15159 15338 15193
rect 15304 15091 15338 15125
rect 15304 15023 15338 15057
rect 15304 14955 15338 14989
rect 15304 14887 15338 14921
rect 15304 14819 15338 14853
rect 15304 14751 15338 14785
rect 15304 14683 15338 14717
rect 15304 14615 15338 14649
rect 15304 14547 15338 14581
rect 15304 14479 15338 14513
rect 15304 14411 15338 14445
rect 15304 14343 15338 14377
rect 15304 14275 15338 14309
rect 15304 14207 15338 14241
rect 15304 14139 15338 14173
rect 15304 14071 15338 14105
rect 15304 14003 15338 14037
rect 15304 13935 15338 13969
rect 15304 13867 15338 13901
rect 14308 13764 14342 13833
rect 14454 13832 14470 13866
rect 14504 13832 14520 13866
rect 14646 13832 14662 13866
rect 14696 13832 14712 13866
rect 14838 13832 14854 13866
rect 14888 13832 14904 13866
rect 15030 13832 15046 13866
rect 15080 13832 15096 13866
rect 15304 13764 15338 13833
rect 14308 13730 14432 13764
rect 14466 13730 14500 13764
rect 14534 13730 14568 13764
rect 14602 13730 14636 13764
rect 14670 13730 14704 13764
rect 14738 13730 14772 13764
rect 14806 13730 14840 13764
rect 14874 13730 14908 13764
rect 14942 13730 14976 13764
rect 15010 13730 15044 13764
rect 15078 13730 15112 13764
rect 15146 13730 15180 13764
rect 15214 13730 15338 13764
rect 16018 16060 16132 16094
rect 16166 16060 16200 16094
rect 16234 16060 16348 16094
rect 16940 16092 17100 16126
rect 17134 16092 17168 16126
rect 17202 16092 17236 16126
rect 17270 16092 17304 16126
rect 17338 16092 17372 16126
rect 17406 16093 17561 16126
rect 17406 16092 17528 16093
rect 16940 16060 17240 16092
rect 16018 15983 16052 16060
rect 16314 15983 16348 16060
rect 16018 15915 16052 15949
rect 16018 15847 16052 15881
rect 16018 15779 16052 15813
rect 16018 15711 16052 15745
rect 16018 15643 16052 15677
rect 16018 15575 16052 15609
rect 16018 15507 16052 15541
rect 16314 15915 16348 15949
rect 16314 15847 16348 15881
rect 16314 15779 16348 15813
rect 16314 15711 16348 15745
rect 16314 15643 16348 15677
rect 16314 15575 16348 15609
rect 16018 15439 16052 15473
rect 16018 15371 16052 15405
rect 16018 15303 16052 15337
rect 16018 15235 16052 15269
rect 16018 15167 16052 15201
rect 16018 15099 16052 15133
rect 16018 15031 16052 15065
rect 16018 14963 16052 14997
rect 16018 14895 16052 14929
rect 16018 14827 16052 14861
rect 16018 14759 16052 14793
rect 16018 14691 16052 14725
rect 16018 14623 16052 14657
rect 16018 14555 16052 14589
rect 16018 14487 16052 14521
rect 16018 14419 16052 14453
rect 16018 14351 16052 14385
rect 16018 14283 16052 14317
rect 16314 15507 16348 15541
rect 16314 15439 16348 15473
rect 16314 15371 16348 15405
rect 16314 15303 16348 15337
rect 16314 15235 16348 15269
rect 16314 15167 16348 15201
rect 16314 15099 16348 15133
rect 16314 15031 16348 15065
rect 16314 14963 16348 14997
rect 16314 14895 16348 14929
rect 16314 14827 16348 14861
rect 16314 14759 16348 14793
rect 16314 14691 16348 14725
rect 16314 14623 16348 14657
rect 16314 14555 16348 14589
rect 16314 14487 16348 14521
rect 16314 14419 16348 14453
rect 16314 14351 16348 14385
rect 16018 14215 16052 14249
rect 16018 14147 16052 14181
rect 16018 14079 16052 14113
rect 16018 14011 16052 14045
rect 16018 13943 16052 13977
rect 16018 13875 16052 13909
rect 16314 14283 16348 14317
rect 16314 14215 16348 14249
rect 16314 14147 16348 14181
rect 16314 14079 16348 14113
rect 16314 14011 16348 14045
rect 16314 13943 16348 13977
rect 16314 13875 16348 13909
rect 16018 13764 16052 13841
rect 16314 13764 16348 13841
rect 16018 13730 16132 13764
rect 16166 13730 16200 13764
rect 16234 13730 16348 13764
rect 16978 16014 17012 16060
rect 17220 15990 17236 16024
rect 17270 15990 17286 16024
rect 17494 16014 17528 16092
rect 16978 15946 17012 15980
rect 16978 15878 17012 15912
rect 16978 15810 17012 15844
rect 16978 15742 17012 15776
rect 16978 15674 17012 15708
rect 16978 15606 17012 15640
rect 16978 15538 17012 15572
rect 16978 15470 17012 15504
rect 16978 15402 17012 15436
rect 16978 15334 17012 15368
rect 16978 15266 17012 15300
rect 16978 15198 17012 15232
rect 16978 15130 17012 15164
rect 16978 15062 17012 15096
rect 16978 14994 17012 15028
rect 16978 14926 17012 14960
rect 16978 14858 17012 14892
rect 16978 14790 17012 14824
rect 16978 14722 17012 14756
rect 16978 14654 17012 14688
rect 16978 14586 17012 14620
rect 16978 14518 17012 14552
rect 16978 14450 17012 14484
rect 16978 14382 17012 14416
rect 16978 14314 17012 14348
rect 16978 14246 17012 14280
rect 16978 14178 17012 14212
rect 16978 14110 17012 14144
rect 16978 14042 17012 14076
rect 16978 13974 17012 14008
rect 16978 13906 17012 13940
rect 17092 15912 17126 15947
rect 17092 15844 17126 15862
rect 17092 15776 17126 15790
rect 17092 15708 17126 15718
rect 17092 15640 17126 15646
rect 17092 15572 17126 15574
rect 17092 15536 17126 15538
rect 17092 15464 17126 15470
rect 17092 15392 17126 15402
rect 17092 15320 17126 15334
rect 17092 15248 17126 15266
rect 17092 15176 17126 15198
rect 17092 15104 17126 15130
rect 17092 15032 17126 15062
rect 17092 14960 17126 14994
rect 17092 14892 17126 14926
rect 17092 14824 17126 14854
rect 17092 14756 17126 14782
rect 17092 14688 17126 14710
rect 17092 14620 17126 14638
rect 17092 14552 17126 14566
rect 17092 14484 17126 14494
rect 17092 14416 17126 14422
rect 17092 14348 17126 14350
rect 17092 14312 17126 14314
rect 17092 14240 17126 14246
rect 17092 14168 17126 14178
rect 17092 14096 17126 14110
rect 17092 14024 17126 14042
rect 17092 13939 17126 13974
rect 17188 15912 17222 15947
rect 17188 15844 17222 15862
rect 17188 15776 17222 15790
rect 17188 15708 17222 15718
rect 17188 15640 17222 15646
rect 17188 15572 17222 15574
rect 17188 15536 17222 15538
rect 17188 15464 17222 15470
rect 17188 15392 17222 15402
rect 17188 15320 17222 15334
rect 17188 15248 17222 15266
rect 17188 15176 17222 15198
rect 17188 15104 17222 15130
rect 17188 15032 17222 15062
rect 17188 14960 17222 14994
rect 17188 14892 17222 14926
rect 17188 14824 17222 14854
rect 17188 14756 17222 14782
rect 17188 14688 17222 14710
rect 17188 14620 17222 14638
rect 17188 14552 17222 14566
rect 17188 14484 17222 14494
rect 17188 14416 17222 14422
rect 17188 14348 17222 14350
rect 17188 14312 17222 14314
rect 17188 14240 17222 14246
rect 17188 14168 17222 14178
rect 17188 14096 17222 14110
rect 17188 14024 17222 14042
rect 17188 13939 17222 13974
rect 17284 15912 17318 15947
rect 17380 15943 17414 15947
rect 17494 15946 17528 15980
rect 17284 15844 17318 15862
rect 17378 15912 17494 15943
rect 17528 15912 17530 15943
rect 17378 15862 17380 15912
rect 17414 15878 17530 15912
rect 17414 15862 17494 15878
rect 17378 15844 17494 15862
rect 17528 15844 17530 15878
rect 17378 15824 17380 15844
rect 17414 15824 17530 15844
rect 17284 15776 17318 15790
rect 17284 15708 17318 15718
rect 17284 15640 17318 15646
rect 17284 15572 17318 15574
rect 17284 15536 17318 15538
rect 17284 15464 17318 15470
rect 17284 15392 17318 15402
rect 17284 15320 17318 15334
rect 17284 15248 17318 15266
rect 17284 15176 17318 15198
rect 17284 15104 17318 15130
rect 17284 15032 17318 15062
rect 17284 14960 17318 14994
rect 17284 14892 17318 14926
rect 17284 14824 17318 14854
rect 17284 14756 17318 14782
rect 17284 14688 17318 14710
rect 17284 14620 17318 14638
rect 17284 14552 17318 14566
rect 17284 14484 17318 14494
rect 17284 14416 17318 14422
rect 17284 14348 17318 14350
rect 17284 14312 17318 14314
rect 17284 14240 17318 14246
rect 17284 14168 17318 14178
rect 17284 14096 17318 14110
rect 17284 14024 17318 14042
rect 17284 13939 17318 13974
rect 17380 15776 17414 15790
rect 17380 15708 17414 15718
rect 17380 15640 17414 15646
rect 17380 15572 17414 15574
rect 17380 15536 17414 15538
rect 17380 15464 17414 15470
rect 17380 15392 17414 15402
rect 17380 15320 17414 15334
rect 17380 15248 17414 15266
rect 17380 15176 17414 15198
rect 17380 15104 17414 15130
rect 17380 15032 17414 15062
rect 17380 14960 17414 14994
rect 17380 14892 17414 14926
rect 17380 14824 17414 14854
rect 17380 14756 17414 14782
rect 17380 14688 17414 14710
rect 17380 14620 17414 14638
rect 17380 14552 17414 14566
rect 17380 14484 17414 14494
rect 17380 14416 17414 14422
rect 17380 14348 17414 14350
rect 17380 14312 17414 14314
rect 17380 14240 17414 14246
rect 17380 14168 17414 14178
rect 17380 14096 17414 14110
rect 17380 14024 17414 14042
rect 17380 13939 17414 13974
rect 17494 15810 17528 15824
rect 17494 15742 17528 15776
rect 17494 15674 17528 15708
rect 17494 15606 17528 15640
rect 17494 15538 17528 15572
rect 17494 15470 17528 15504
rect 17494 15402 17528 15436
rect 17494 15334 17528 15368
rect 17494 15266 17528 15300
rect 17494 15198 17528 15232
rect 17494 15130 17528 15164
rect 17494 15062 17528 15096
rect 17494 14994 17528 15028
rect 17494 14926 17528 14960
rect 17494 14858 17528 14892
rect 17494 14790 17528 14824
rect 17494 14722 17528 14756
rect 17494 14654 17528 14688
rect 17494 14586 17528 14620
rect 17494 14518 17528 14552
rect 17494 14450 17528 14484
rect 17494 14382 17528 14416
rect 17494 14314 17528 14348
rect 17494 14246 17528 14280
rect 17494 14178 17528 14212
rect 17494 14110 17528 14144
rect 17494 14042 17528 14076
rect 17494 13974 17528 14008
rect 17494 13906 17528 13940
rect 16978 13794 17012 13872
rect 17124 13862 17140 13896
rect 17174 13862 17190 13896
rect 17316 13862 17332 13896
rect 17366 13862 17382 13896
rect 17494 13794 17528 13872
rect 16978 13760 17100 13794
rect 17134 13760 17168 13794
rect 17202 13760 17236 13794
rect 17270 13760 17304 13794
rect 17338 13760 17372 13794
rect 17406 13760 17528 13794
rect 13074 13546 17870 13590
rect 13074 13512 13329 13546
rect 13363 13512 13397 13546
rect 13431 13512 13465 13546
rect 13499 13512 13533 13546
rect 13567 13512 13601 13546
rect 13635 13512 13669 13546
rect 13703 13512 13737 13546
rect 13771 13512 13805 13546
rect 13839 13512 13873 13546
rect 13907 13512 13941 13546
rect 13975 13512 14009 13546
rect 14043 13512 14077 13546
rect 14111 13512 14145 13546
rect 14179 13512 14213 13546
rect 14247 13512 14281 13546
rect 14315 13512 14349 13546
rect 14383 13512 14417 13546
rect 14451 13512 14485 13546
rect 14519 13512 14553 13546
rect 14587 13512 14621 13546
rect 14655 13512 14689 13546
rect 14723 13512 14757 13546
rect 14791 13512 14825 13546
rect 14859 13512 14893 13546
rect 14927 13512 14961 13546
rect 14995 13512 15029 13546
rect 15063 13512 15097 13546
rect 15131 13512 15165 13546
rect 15199 13512 15233 13546
rect 15267 13512 15301 13546
rect 15335 13512 15369 13546
rect 15403 13512 15437 13546
rect 15471 13512 15505 13546
rect 15539 13512 15573 13546
rect 15607 13512 15641 13546
rect 15675 13512 15709 13546
rect 15743 13512 15777 13546
rect 15811 13512 15845 13546
rect 15879 13512 15913 13546
rect 15947 13512 15981 13546
rect 16015 13512 16049 13546
rect 16083 13512 16117 13546
rect 16151 13512 16185 13546
rect 16219 13512 16253 13546
rect 16287 13512 16321 13546
rect 16355 13512 16389 13546
rect 16423 13512 16457 13546
rect 16491 13512 16525 13546
rect 16559 13512 16593 13546
rect 16627 13512 16661 13546
rect 16695 13512 16729 13546
rect 16763 13512 16797 13546
rect 16831 13512 16865 13546
rect 16899 13512 16933 13546
rect 16967 13512 17001 13546
rect 17035 13512 17069 13546
rect 17103 13512 17137 13546
rect 17171 13512 17205 13546
rect 17239 13512 17273 13546
rect 17307 13512 17341 13546
rect 17375 13512 17409 13546
rect 17443 13512 17477 13546
rect 17511 13512 17545 13546
rect 17579 13512 17870 13546
rect 13074 13455 17870 13512
rect 13074 13416 13209 13455
rect 13074 13382 13122 13416
rect 13156 13382 13209 13416
rect 13074 13348 13209 13382
rect 17728 13425 17870 13455
rect 17728 13391 17785 13425
rect 17819 13391 17870 13425
rect 17728 13357 17870 13391
rect 13074 13314 13122 13348
rect 13156 13314 13209 13348
rect 13074 13280 13209 13314
rect 13074 13246 13122 13280
rect 13156 13246 13209 13280
rect 13074 13212 13209 13246
rect 16122 13331 16242 13354
rect 16122 13297 16165 13331
rect 16199 13297 16242 13331
rect 13074 13178 13122 13212
rect 13156 13178 13209 13212
rect 13074 13144 13209 13178
rect 13074 13110 13122 13144
rect 13156 13110 13209 13144
rect 13480 13181 13571 13215
rect 16122 13198 16242 13297
rect 17000 13310 17118 13334
rect 17000 13276 17040 13310
rect 17074 13276 17118 13310
rect 17000 13254 17118 13276
rect 17728 13323 17785 13357
rect 17819 13323 17870 13357
rect 17728 13289 17870 13323
rect 17728 13255 17785 13289
rect 17819 13255 17870 13289
rect 17728 13221 17870 13255
rect 13480 13147 13509 13181
rect 13543 13147 13571 13181
rect 13480 13115 13571 13147
rect 13614 13171 17474 13198
rect 13614 13137 13695 13171
rect 13729 13167 17474 13171
rect 13729 13137 14049 13167
rect 13614 13133 14049 13137
rect 14083 13166 15460 13167
rect 14083 13165 14755 13166
rect 14083 13133 14402 13165
rect 13614 13131 14402 13133
rect 14436 13132 14755 13165
rect 14789 13132 15106 13166
rect 15140 13133 15460 13166
rect 15494 13166 17474 13167
rect 15494 13133 15810 13166
rect 15140 13132 15810 13133
rect 15844 13165 17474 13166
rect 15844 13132 16162 13165
rect 14436 13131 16162 13132
rect 16196 13131 16515 13165
rect 16549 13131 16864 13165
rect 16898 13131 17218 13165
rect 17252 13131 17391 13165
rect 17425 13131 17474 13165
rect 13614 13119 17474 13131
rect 17728 13187 17785 13221
rect 17819 13187 17870 13221
rect 17728 13153 17870 13187
rect 17728 13119 17785 13153
rect 17819 13119 17870 13153
rect 13675 13115 13750 13119
rect 14029 13111 14104 13119
rect 13074 13076 13209 13110
rect 14382 13109 14457 13119
rect 14735 13110 14810 13119
rect 15086 13110 15161 13119
rect 15440 13111 15515 13119
rect 15790 13110 15865 13119
rect 16122 13114 16242 13119
rect 16142 13109 16217 13114
rect 16495 13109 16570 13119
rect 16844 13109 16919 13119
rect 17198 13109 17273 13119
rect 17371 13109 17446 13119
rect 13074 13042 13122 13076
rect 13156 13042 13209 13076
rect 17728 13085 17870 13119
rect 13074 13008 13209 13042
rect 13074 12974 13122 13008
rect 13156 12974 13209 13008
rect 13074 12940 13209 12974
rect 13074 12906 13122 12940
rect 13156 12906 13209 12940
rect 13074 12872 13209 12906
rect 13074 12838 13122 12872
rect 13156 12838 13209 12872
rect 13074 12804 13209 12838
rect 13074 12770 13122 12804
rect 13156 12770 13209 12804
rect 13074 12736 13209 12770
rect 13074 12702 13122 12736
rect 13156 12702 13209 12736
rect 13074 12668 13209 12702
rect 13074 12634 13122 12668
rect 13156 12634 13209 12668
rect 13074 12600 13209 12634
rect 13074 12566 13122 12600
rect 13156 12566 13209 12600
rect 13074 12532 13209 12566
rect 13074 12498 13122 12532
rect 13156 12498 13209 12532
rect 13074 12464 13209 12498
rect 13074 12430 13122 12464
rect 13156 12430 13209 12464
rect 13074 12396 13209 12430
rect 13074 12362 13122 12396
rect 13156 12362 13209 12396
rect 13074 12328 13209 12362
rect 13074 12294 13122 12328
rect 13156 12294 13209 12328
rect 13074 12260 13209 12294
rect 13074 12226 13122 12260
rect 13156 12226 13209 12260
rect 13074 12192 13209 12226
rect 13074 12158 13122 12192
rect 13156 12158 13209 12192
rect 13074 12124 13209 12158
rect 13074 12090 13122 12124
rect 13156 12090 13209 12124
rect 13074 12056 13209 12090
rect 13074 12022 13122 12056
rect 13156 12022 13209 12056
rect 13074 11988 13209 12022
rect 13074 11954 13122 11988
rect 13156 11954 13209 11988
rect 13074 11920 13209 11954
rect 13074 11886 13122 11920
rect 13156 11886 13209 11920
rect 13074 11852 13209 11886
rect 13074 11818 13122 11852
rect 13156 11818 13209 11852
rect 13074 11784 13209 11818
rect 13074 11750 13122 11784
rect 13156 11750 13209 11784
rect 13074 11716 13209 11750
rect 13074 11682 13122 11716
rect 13156 11682 13209 11716
rect 13074 11648 13209 11682
rect 13074 11614 13122 11648
rect 13156 11614 13209 11648
rect 13074 11580 13209 11614
rect 13074 11546 13122 11580
rect 13156 11546 13209 11580
rect 13074 11512 13209 11546
rect 13074 11478 13122 11512
rect 13156 11478 13209 11512
rect 13074 11444 13209 11478
rect 13074 11410 13122 11444
rect 13156 11410 13209 11444
rect 13074 11376 13209 11410
rect 13074 11342 13122 11376
rect 13156 11342 13209 11376
rect 13074 11308 13209 11342
rect 13074 11274 13122 11308
rect 13156 11274 13209 11308
rect 13074 11240 13209 11274
rect 13074 11206 13122 11240
rect 13156 11206 13209 11240
rect 13074 11172 13209 11206
rect 13074 11138 13122 11172
rect 13156 11138 13209 11172
rect 13074 11104 13209 11138
rect 13074 11070 13122 11104
rect 13156 11070 13209 11104
rect 13074 11036 13209 11070
rect 13434 13039 13468 13074
rect 13434 12971 13468 12989
rect 13434 12903 13468 12917
rect 13434 12835 13468 12845
rect 13434 12767 13468 12773
rect 13434 12699 13468 12701
rect 13434 12663 13468 12665
rect 13434 12591 13468 12597
rect 13434 12519 13468 12529
rect 13434 12447 13468 12461
rect 13434 12375 13468 12393
rect 13434 12303 13468 12325
rect 13434 12231 13468 12257
rect 13434 12159 13468 12189
rect 13434 12087 13468 12121
rect 13434 12019 13468 12053
rect 13434 11951 13468 11981
rect 13434 11883 13468 11909
rect 13434 11815 13468 11837
rect 13434 11747 13468 11765
rect 13434 11679 13468 11693
rect 13434 11611 13468 11621
rect 13434 11543 13468 11549
rect 13434 11475 13468 11477
rect 13434 11439 13468 11441
rect 13434 11367 13468 11373
rect 13434 11295 13468 11305
rect 13434 11223 13468 11237
rect 13434 11151 13468 11169
rect 13434 11066 13468 11101
rect 13522 13039 13556 13074
rect 13522 12971 13556 12989
rect 13522 12903 13556 12917
rect 13522 12835 13556 12845
rect 13522 12767 13556 12773
rect 13522 12699 13556 12701
rect 13522 12663 13556 12665
rect 13522 12591 13556 12597
rect 13522 12519 13556 12529
rect 13522 12447 13556 12461
rect 13522 12375 13556 12393
rect 13522 12303 13556 12325
rect 13522 12231 13556 12257
rect 13522 12159 13556 12189
rect 13522 12087 13556 12121
rect 13522 12019 13556 12053
rect 13522 11951 13556 11981
rect 13522 11883 13556 11909
rect 13522 11815 13556 11837
rect 13522 11747 13556 11765
rect 13522 11679 13556 11693
rect 13522 11611 13556 11621
rect 13522 11543 13556 11549
rect 13522 11475 13556 11477
rect 13522 11439 13556 11441
rect 13522 11367 13556 11373
rect 13522 11295 13556 11305
rect 13522 11223 13556 11237
rect 13522 11151 13556 11169
rect 13522 11066 13556 11101
rect 13610 13039 13644 13074
rect 13610 12971 13644 12989
rect 13610 12903 13644 12917
rect 13610 12835 13644 12845
rect 13610 12767 13644 12773
rect 13610 12699 13644 12701
rect 13610 12663 13644 12665
rect 13610 12591 13644 12597
rect 13610 12519 13644 12529
rect 13610 12447 13644 12461
rect 13610 12375 13644 12393
rect 13610 12303 13644 12325
rect 13610 12231 13644 12257
rect 13610 12159 13644 12189
rect 13610 12087 13644 12121
rect 13610 12019 13644 12053
rect 13610 11951 13644 11981
rect 13610 11883 13644 11909
rect 13610 11815 13644 11837
rect 13610 11747 13644 11765
rect 13610 11679 13644 11693
rect 13610 11611 13644 11621
rect 13610 11543 13644 11549
rect 13610 11475 13644 11477
rect 13610 11439 13644 11441
rect 13610 11367 13644 11373
rect 13610 11295 13644 11305
rect 13610 11223 13644 11237
rect 13610 11151 13644 11169
rect 13610 11066 13644 11101
rect 13698 13039 13732 13074
rect 13698 12971 13732 12989
rect 13698 12903 13732 12917
rect 13698 12835 13732 12845
rect 13698 12767 13732 12773
rect 13698 12699 13732 12701
rect 13698 12663 13732 12665
rect 13698 12591 13732 12597
rect 13698 12519 13732 12529
rect 13698 12447 13732 12461
rect 13698 12375 13732 12393
rect 13698 12303 13732 12325
rect 13698 12231 13732 12257
rect 13698 12159 13732 12189
rect 13698 12087 13732 12121
rect 13698 12019 13732 12053
rect 13698 11951 13732 11981
rect 13698 11883 13732 11909
rect 13698 11815 13732 11837
rect 13698 11747 13732 11765
rect 13698 11679 13732 11693
rect 13698 11611 13732 11621
rect 13698 11543 13732 11549
rect 13698 11475 13732 11477
rect 13698 11439 13732 11441
rect 13698 11367 13732 11373
rect 13698 11295 13732 11305
rect 13698 11223 13732 11237
rect 13698 11151 13732 11169
rect 13698 11066 13732 11101
rect 13786 13039 13820 13074
rect 13786 12971 13820 12989
rect 13786 12903 13820 12917
rect 13786 12835 13820 12845
rect 13786 12767 13820 12773
rect 13786 12699 13820 12701
rect 13786 12663 13820 12665
rect 13786 12591 13820 12597
rect 13786 12519 13820 12529
rect 13786 12447 13820 12461
rect 13786 12375 13820 12393
rect 13786 12303 13820 12325
rect 13786 12231 13820 12257
rect 13786 12159 13820 12189
rect 13786 12087 13820 12121
rect 13786 12019 13820 12053
rect 13786 11951 13820 11981
rect 13786 11883 13820 11909
rect 13786 11815 13820 11837
rect 13786 11747 13820 11765
rect 13786 11679 13820 11693
rect 13786 11611 13820 11621
rect 13786 11543 13820 11549
rect 13786 11475 13820 11477
rect 13786 11439 13820 11441
rect 13786 11367 13820 11373
rect 13786 11295 13820 11305
rect 13786 11223 13820 11237
rect 13786 11151 13820 11169
rect 13786 11066 13820 11101
rect 13874 13039 13908 13074
rect 13874 12971 13908 12989
rect 13874 12903 13908 12917
rect 13874 12835 13908 12845
rect 13874 12767 13908 12773
rect 13874 12699 13908 12701
rect 13874 12663 13908 12665
rect 13874 12591 13908 12597
rect 13874 12519 13908 12529
rect 13874 12447 13908 12461
rect 13874 12375 13908 12393
rect 13874 12303 13908 12325
rect 13874 12231 13908 12257
rect 13874 12159 13908 12189
rect 13874 12087 13908 12121
rect 13874 12019 13908 12053
rect 13874 11951 13908 11981
rect 13874 11883 13908 11909
rect 13874 11815 13908 11837
rect 13874 11747 13908 11765
rect 13874 11679 13908 11693
rect 13874 11611 13908 11621
rect 13874 11543 13908 11549
rect 13874 11475 13908 11477
rect 13874 11439 13908 11441
rect 13874 11367 13908 11373
rect 13874 11295 13908 11305
rect 13874 11223 13908 11237
rect 13874 11151 13908 11169
rect 13874 11066 13908 11101
rect 13962 13039 13996 13074
rect 13962 12971 13996 12989
rect 13962 12903 13996 12917
rect 13962 12835 13996 12845
rect 13962 12767 13996 12773
rect 13962 12699 13996 12701
rect 13962 12663 13996 12665
rect 13962 12591 13996 12597
rect 13962 12519 13996 12529
rect 13962 12447 13996 12461
rect 13962 12375 13996 12393
rect 13962 12303 13996 12325
rect 13962 12231 13996 12257
rect 13962 12159 13996 12189
rect 13962 12087 13996 12121
rect 13962 12019 13996 12053
rect 13962 11951 13996 11981
rect 13962 11883 13996 11909
rect 13962 11815 13996 11837
rect 13962 11747 13996 11765
rect 13962 11679 13996 11693
rect 13962 11611 13996 11621
rect 13962 11543 13996 11549
rect 13962 11475 13996 11477
rect 13962 11439 13996 11441
rect 13962 11367 13996 11373
rect 13962 11295 13996 11305
rect 13962 11223 13996 11237
rect 13962 11151 13996 11169
rect 13962 11066 13996 11101
rect 14050 13039 14084 13074
rect 14050 12971 14084 12989
rect 14050 12903 14084 12917
rect 14050 12835 14084 12845
rect 14050 12767 14084 12773
rect 14050 12699 14084 12701
rect 14050 12663 14084 12665
rect 14050 12591 14084 12597
rect 14050 12519 14084 12529
rect 14050 12447 14084 12461
rect 14050 12375 14084 12393
rect 14050 12303 14084 12325
rect 14050 12231 14084 12257
rect 14050 12159 14084 12189
rect 14050 12087 14084 12121
rect 14050 12019 14084 12053
rect 14050 11951 14084 11981
rect 14050 11883 14084 11909
rect 14050 11815 14084 11837
rect 14050 11747 14084 11765
rect 14050 11679 14084 11693
rect 14050 11611 14084 11621
rect 14050 11543 14084 11549
rect 14050 11475 14084 11477
rect 14050 11439 14084 11441
rect 14050 11367 14084 11373
rect 14050 11295 14084 11305
rect 14050 11223 14084 11237
rect 14050 11151 14084 11169
rect 14050 11066 14084 11101
rect 14138 13039 14172 13074
rect 14138 12971 14172 12989
rect 14138 12903 14172 12917
rect 14138 12835 14172 12845
rect 14138 12767 14172 12773
rect 14138 12699 14172 12701
rect 14138 12663 14172 12665
rect 14138 12591 14172 12597
rect 14138 12519 14172 12529
rect 14138 12447 14172 12461
rect 14138 12375 14172 12393
rect 14138 12303 14172 12325
rect 14138 12231 14172 12257
rect 14138 12159 14172 12189
rect 14138 12087 14172 12121
rect 14138 12019 14172 12053
rect 14138 11951 14172 11981
rect 14138 11883 14172 11909
rect 14138 11815 14172 11837
rect 14138 11747 14172 11765
rect 14138 11679 14172 11693
rect 14138 11611 14172 11621
rect 14138 11543 14172 11549
rect 14138 11475 14172 11477
rect 14138 11439 14172 11441
rect 14138 11367 14172 11373
rect 14138 11295 14172 11305
rect 14138 11223 14172 11237
rect 14138 11151 14172 11169
rect 14138 11066 14172 11101
rect 14226 13039 14260 13074
rect 14226 12971 14260 12989
rect 14226 12903 14260 12917
rect 14226 12835 14260 12845
rect 14226 12767 14260 12773
rect 14226 12699 14260 12701
rect 14226 12663 14260 12665
rect 14226 12591 14260 12597
rect 14226 12519 14260 12529
rect 14226 12447 14260 12461
rect 14226 12375 14260 12393
rect 14226 12303 14260 12325
rect 14226 12231 14260 12257
rect 14226 12159 14260 12189
rect 14226 12087 14260 12121
rect 14226 12019 14260 12053
rect 14226 11951 14260 11981
rect 14226 11883 14260 11909
rect 14226 11815 14260 11837
rect 14226 11747 14260 11765
rect 14226 11679 14260 11693
rect 14226 11611 14260 11621
rect 14226 11543 14260 11549
rect 14226 11475 14260 11477
rect 14226 11439 14260 11441
rect 14226 11367 14260 11373
rect 14226 11295 14260 11305
rect 14226 11223 14260 11237
rect 14226 11151 14260 11169
rect 14226 11066 14260 11101
rect 14314 13039 14348 13074
rect 14314 12971 14348 12989
rect 14314 12903 14348 12917
rect 14314 12835 14348 12845
rect 14314 12767 14348 12773
rect 14314 12699 14348 12701
rect 14314 12663 14348 12665
rect 14314 12591 14348 12597
rect 14314 12519 14348 12529
rect 14314 12447 14348 12461
rect 14314 12375 14348 12393
rect 14314 12303 14348 12325
rect 14314 12231 14348 12257
rect 14314 12159 14348 12189
rect 14314 12087 14348 12121
rect 14314 12019 14348 12053
rect 14314 11951 14348 11981
rect 14314 11883 14348 11909
rect 14314 11815 14348 11837
rect 14314 11747 14348 11765
rect 14314 11679 14348 11693
rect 14314 11611 14348 11621
rect 14314 11543 14348 11549
rect 14314 11475 14348 11477
rect 14314 11439 14348 11441
rect 14314 11367 14348 11373
rect 14314 11295 14348 11305
rect 14314 11223 14348 11237
rect 14314 11151 14348 11169
rect 14314 11066 14348 11101
rect 14402 13039 14436 13074
rect 14402 12971 14436 12989
rect 14402 12903 14436 12917
rect 14402 12835 14436 12845
rect 14402 12767 14436 12773
rect 14402 12699 14436 12701
rect 14402 12663 14436 12665
rect 14402 12591 14436 12597
rect 14402 12519 14436 12529
rect 14402 12447 14436 12461
rect 14402 12375 14436 12393
rect 14402 12303 14436 12325
rect 14402 12231 14436 12257
rect 14402 12159 14436 12189
rect 14402 12087 14436 12121
rect 14402 12019 14436 12053
rect 14402 11951 14436 11981
rect 14402 11883 14436 11909
rect 14402 11815 14436 11837
rect 14402 11747 14436 11765
rect 14402 11679 14436 11693
rect 14402 11611 14436 11621
rect 14402 11543 14436 11549
rect 14402 11475 14436 11477
rect 14402 11439 14436 11441
rect 14402 11367 14436 11373
rect 14402 11295 14436 11305
rect 14402 11223 14436 11237
rect 14402 11151 14436 11169
rect 14402 11066 14436 11101
rect 14490 13039 14524 13074
rect 14490 12971 14524 12989
rect 14490 12903 14524 12917
rect 14490 12835 14524 12845
rect 14490 12767 14524 12773
rect 14490 12699 14524 12701
rect 14490 12663 14524 12665
rect 14490 12591 14524 12597
rect 14490 12519 14524 12529
rect 14490 12447 14524 12461
rect 14490 12375 14524 12393
rect 14490 12303 14524 12325
rect 14490 12231 14524 12257
rect 14490 12159 14524 12189
rect 14490 12087 14524 12121
rect 14490 12019 14524 12053
rect 14490 11951 14524 11981
rect 14490 11883 14524 11909
rect 14490 11815 14524 11837
rect 14490 11747 14524 11765
rect 14490 11679 14524 11693
rect 14490 11611 14524 11621
rect 14490 11543 14524 11549
rect 14490 11475 14524 11477
rect 14490 11439 14524 11441
rect 14490 11367 14524 11373
rect 14490 11295 14524 11305
rect 14490 11223 14524 11237
rect 14490 11151 14524 11169
rect 14490 11066 14524 11101
rect 14578 13039 14612 13074
rect 14578 12971 14612 12989
rect 14578 12903 14612 12917
rect 14578 12835 14612 12845
rect 14578 12767 14612 12773
rect 14578 12699 14612 12701
rect 14578 12663 14612 12665
rect 14578 12591 14612 12597
rect 14578 12519 14612 12529
rect 14578 12447 14612 12461
rect 14578 12375 14612 12393
rect 14578 12303 14612 12325
rect 14578 12231 14612 12257
rect 14578 12159 14612 12189
rect 14578 12087 14612 12121
rect 14578 12019 14612 12053
rect 14578 11951 14612 11981
rect 14578 11883 14612 11909
rect 14578 11815 14612 11837
rect 14578 11747 14612 11765
rect 14578 11679 14612 11693
rect 14578 11611 14612 11621
rect 14578 11543 14612 11549
rect 14578 11475 14612 11477
rect 14578 11439 14612 11441
rect 14578 11367 14612 11373
rect 14578 11295 14612 11305
rect 14578 11223 14612 11237
rect 14578 11151 14612 11169
rect 14578 11066 14612 11101
rect 14666 13039 14700 13074
rect 14666 12971 14700 12989
rect 14666 12903 14700 12917
rect 14666 12835 14700 12845
rect 14666 12767 14700 12773
rect 14666 12699 14700 12701
rect 14666 12663 14700 12665
rect 14666 12591 14700 12597
rect 14666 12519 14700 12529
rect 14666 12447 14700 12461
rect 14666 12375 14700 12393
rect 14666 12303 14700 12325
rect 14666 12231 14700 12257
rect 14666 12159 14700 12189
rect 14666 12087 14700 12121
rect 14666 12019 14700 12053
rect 14666 11951 14700 11981
rect 14666 11883 14700 11909
rect 14666 11815 14700 11837
rect 14666 11747 14700 11765
rect 14666 11679 14700 11693
rect 14666 11611 14700 11621
rect 14666 11543 14700 11549
rect 14666 11475 14700 11477
rect 14666 11439 14700 11441
rect 14666 11367 14700 11373
rect 14666 11295 14700 11305
rect 14666 11223 14700 11237
rect 14666 11151 14700 11169
rect 14666 11066 14700 11101
rect 14754 13039 14788 13074
rect 14754 12971 14788 12989
rect 14754 12903 14788 12917
rect 14754 12835 14788 12845
rect 14754 12767 14788 12773
rect 14754 12699 14788 12701
rect 14754 12663 14788 12665
rect 14754 12591 14788 12597
rect 14754 12519 14788 12529
rect 14754 12447 14788 12461
rect 14754 12375 14788 12393
rect 14754 12303 14788 12325
rect 14754 12231 14788 12257
rect 14754 12159 14788 12189
rect 14754 12087 14788 12121
rect 14754 12019 14788 12053
rect 14754 11951 14788 11981
rect 14754 11883 14788 11909
rect 14754 11815 14788 11837
rect 14754 11747 14788 11765
rect 14754 11679 14788 11693
rect 14754 11611 14788 11621
rect 14754 11543 14788 11549
rect 14754 11475 14788 11477
rect 14754 11439 14788 11441
rect 14754 11367 14788 11373
rect 14754 11295 14788 11305
rect 14754 11223 14788 11237
rect 14754 11151 14788 11169
rect 14754 11066 14788 11101
rect 14842 13039 14876 13074
rect 14842 12971 14876 12989
rect 14842 12903 14876 12917
rect 14842 12835 14876 12845
rect 14842 12767 14876 12773
rect 14842 12699 14876 12701
rect 14842 12663 14876 12665
rect 14842 12591 14876 12597
rect 14842 12519 14876 12529
rect 14842 12447 14876 12461
rect 14842 12375 14876 12393
rect 14842 12303 14876 12325
rect 14842 12231 14876 12257
rect 14842 12159 14876 12189
rect 14842 12087 14876 12121
rect 14842 12019 14876 12053
rect 14842 11951 14876 11981
rect 14842 11883 14876 11909
rect 14842 11815 14876 11837
rect 14842 11747 14876 11765
rect 14842 11679 14876 11693
rect 14842 11611 14876 11621
rect 14842 11543 14876 11549
rect 14842 11475 14876 11477
rect 14842 11439 14876 11441
rect 14842 11367 14876 11373
rect 14842 11295 14876 11305
rect 14842 11223 14876 11237
rect 14842 11151 14876 11169
rect 14842 11066 14876 11101
rect 14930 13039 14964 13074
rect 14930 12971 14964 12989
rect 14930 12903 14964 12917
rect 14930 12835 14964 12845
rect 14930 12767 14964 12773
rect 14930 12699 14964 12701
rect 14930 12663 14964 12665
rect 14930 12591 14964 12597
rect 14930 12519 14964 12529
rect 14930 12447 14964 12461
rect 14930 12375 14964 12393
rect 14930 12303 14964 12325
rect 14930 12231 14964 12257
rect 14930 12159 14964 12189
rect 14930 12087 14964 12121
rect 14930 12019 14964 12053
rect 14930 11951 14964 11981
rect 14930 11883 14964 11909
rect 14930 11815 14964 11837
rect 14930 11747 14964 11765
rect 14930 11679 14964 11693
rect 14930 11611 14964 11621
rect 14930 11543 14964 11549
rect 14930 11475 14964 11477
rect 14930 11439 14964 11441
rect 14930 11367 14964 11373
rect 14930 11295 14964 11305
rect 14930 11223 14964 11237
rect 14930 11151 14964 11169
rect 14930 11066 14964 11101
rect 15018 13039 15052 13074
rect 15018 12971 15052 12989
rect 15018 12903 15052 12917
rect 15018 12835 15052 12845
rect 15018 12767 15052 12773
rect 15018 12699 15052 12701
rect 15018 12663 15052 12665
rect 15018 12591 15052 12597
rect 15018 12519 15052 12529
rect 15018 12447 15052 12461
rect 15018 12375 15052 12393
rect 15018 12303 15052 12325
rect 15018 12231 15052 12257
rect 15018 12159 15052 12189
rect 15018 12087 15052 12121
rect 15018 12019 15052 12053
rect 15018 11951 15052 11981
rect 15018 11883 15052 11909
rect 15018 11815 15052 11837
rect 15018 11747 15052 11765
rect 15018 11679 15052 11693
rect 15018 11611 15052 11621
rect 15018 11543 15052 11549
rect 15018 11475 15052 11477
rect 15018 11439 15052 11441
rect 15018 11367 15052 11373
rect 15018 11295 15052 11305
rect 15018 11223 15052 11237
rect 15018 11151 15052 11169
rect 15018 11066 15052 11101
rect 15106 13039 15140 13074
rect 15106 12971 15140 12989
rect 15106 12903 15140 12917
rect 15106 12835 15140 12845
rect 15106 12767 15140 12773
rect 15106 12699 15140 12701
rect 15106 12663 15140 12665
rect 15106 12591 15140 12597
rect 15106 12519 15140 12529
rect 15106 12447 15140 12461
rect 15106 12375 15140 12393
rect 15106 12303 15140 12325
rect 15106 12231 15140 12257
rect 15106 12159 15140 12189
rect 15106 12087 15140 12121
rect 15106 12019 15140 12053
rect 15106 11951 15140 11981
rect 15106 11883 15140 11909
rect 15106 11815 15140 11837
rect 15106 11747 15140 11765
rect 15106 11679 15140 11693
rect 15106 11611 15140 11621
rect 15106 11543 15140 11549
rect 15106 11475 15140 11477
rect 15106 11439 15140 11441
rect 15106 11367 15140 11373
rect 15106 11295 15140 11305
rect 15106 11223 15140 11237
rect 15106 11151 15140 11169
rect 15106 11066 15140 11101
rect 15194 13039 15228 13074
rect 15194 12971 15228 12989
rect 15194 12903 15228 12917
rect 15194 12835 15228 12845
rect 15194 12767 15228 12773
rect 15194 12699 15228 12701
rect 15194 12663 15228 12665
rect 15194 12591 15228 12597
rect 15194 12519 15228 12529
rect 15194 12447 15228 12461
rect 15194 12375 15228 12393
rect 15194 12303 15228 12325
rect 15194 12231 15228 12257
rect 15194 12159 15228 12189
rect 15194 12087 15228 12121
rect 15194 12019 15228 12053
rect 15194 11951 15228 11981
rect 15194 11883 15228 11909
rect 15194 11815 15228 11837
rect 15194 11747 15228 11765
rect 15194 11679 15228 11693
rect 15194 11611 15228 11621
rect 15194 11543 15228 11549
rect 15194 11475 15228 11477
rect 15194 11439 15228 11441
rect 15194 11367 15228 11373
rect 15194 11295 15228 11305
rect 15194 11223 15228 11237
rect 15194 11151 15228 11169
rect 15194 11066 15228 11101
rect 15282 13039 15316 13074
rect 15282 12971 15316 12989
rect 15282 12903 15316 12917
rect 15282 12835 15316 12845
rect 15282 12767 15316 12773
rect 15282 12699 15316 12701
rect 15282 12663 15316 12665
rect 15282 12591 15316 12597
rect 15282 12519 15316 12529
rect 15282 12447 15316 12461
rect 15282 12375 15316 12393
rect 15282 12303 15316 12325
rect 15282 12231 15316 12257
rect 15282 12159 15316 12189
rect 15282 12087 15316 12121
rect 15282 12019 15316 12053
rect 15282 11951 15316 11981
rect 15282 11883 15316 11909
rect 15282 11815 15316 11837
rect 15282 11747 15316 11765
rect 15282 11679 15316 11693
rect 15282 11611 15316 11621
rect 15282 11543 15316 11549
rect 15282 11475 15316 11477
rect 15282 11439 15316 11441
rect 15282 11367 15316 11373
rect 15282 11295 15316 11305
rect 15282 11223 15316 11237
rect 15282 11151 15316 11169
rect 15282 11066 15316 11101
rect 15370 13039 15404 13074
rect 15370 12971 15404 12989
rect 15370 12903 15404 12917
rect 15370 12835 15404 12845
rect 15370 12767 15404 12773
rect 15370 12699 15404 12701
rect 15370 12663 15404 12665
rect 15370 12591 15404 12597
rect 15370 12519 15404 12529
rect 15370 12447 15404 12461
rect 15370 12375 15404 12393
rect 15370 12303 15404 12325
rect 15370 12231 15404 12257
rect 15370 12159 15404 12189
rect 15370 12087 15404 12121
rect 15370 12019 15404 12053
rect 15370 11951 15404 11981
rect 15370 11883 15404 11909
rect 15370 11815 15404 11837
rect 15370 11747 15404 11765
rect 15370 11679 15404 11693
rect 15370 11611 15404 11621
rect 15370 11543 15404 11549
rect 15370 11475 15404 11477
rect 15370 11439 15404 11441
rect 15370 11367 15404 11373
rect 15370 11295 15404 11305
rect 15370 11223 15404 11237
rect 15370 11151 15404 11169
rect 15370 11066 15404 11101
rect 15458 13039 15492 13074
rect 15458 12971 15492 12989
rect 15458 12903 15492 12917
rect 15458 12835 15492 12845
rect 15458 12767 15492 12773
rect 15458 12699 15492 12701
rect 15458 12663 15492 12665
rect 15458 12591 15492 12597
rect 15458 12519 15492 12529
rect 15458 12447 15492 12461
rect 15458 12375 15492 12393
rect 15458 12303 15492 12325
rect 15458 12231 15492 12257
rect 15458 12159 15492 12189
rect 15458 12087 15492 12121
rect 15458 12019 15492 12053
rect 15458 11951 15492 11981
rect 15458 11883 15492 11909
rect 15458 11815 15492 11837
rect 15458 11747 15492 11765
rect 15458 11679 15492 11693
rect 15458 11611 15492 11621
rect 15458 11543 15492 11549
rect 15458 11475 15492 11477
rect 15458 11439 15492 11441
rect 15458 11367 15492 11373
rect 15458 11295 15492 11305
rect 15458 11223 15492 11237
rect 15458 11151 15492 11169
rect 15458 11066 15492 11101
rect 15546 13039 15580 13074
rect 15546 12971 15580 12989
rect 15546 12903 15580 12917
rect 15546 12835 15580 12845
rect 15546 12767 15580 12773
rect 15546 12699 15580 12701
rect 15546 12663 15580 12665
rect 15546 12591 15580 12597
rect 15546 12519 15580 12529
rect 15546 12447 15580 12461
rect 15546 12375 15580 12393
rect 15546 12303 15580 12325
rect 15546 12231 15580 12257
rect 15546 12159 15580 12189
rect 15546 12087 15580 12121
rect 15546 12019 15580 12053
rect 15546 11951 15580 11981
rect 15546 11883 15580 11909
rect 15546 11815 15580 11837
rect 15546 11747 15580 11765
rect 15546 11679 15580 11693
rect 15546 11611 15580 11621
rect 15546 11543 15580 11549
rect 15546 11475 15580 11477
rect 15546 11439 15580 11441
rect 15546 11367 15580 11373
rect 15546 11295 15580 11305
rect 15546 11223 15580 11237
rect 15546 11151 15580 11169
rect 15546 11066 15580 11101
rect 15634 13039 15668 13074
rect 15634 12971 15668 12989
rect 15634 12903 15668 12917
rect 15634 12835 15668 12845
rect 15634 12767 15668 12773
rect 15634 12699 15668 12701
rect 15634 12663 15668 12665
rect 15634 12591 15668 12597
rect 15634 12519 15668 12529
rect 15634 12447 15668 12461
rect 15634 12375 15668 12393
rect 15634 12303 15668 12325
rect 15634 12231 15668 12257
rect 15634 12159 15668 12189
rect 15634 12087 15668 12121
rect 15634 12019 15668 12053
rect 15634 11951 15668 11981
rect 15634 11883 15668 11909
rect 15634 11815 15668 11837
rect 15634 11747 15668 11765
rect 15634 11679 15668 11693
rect 15634 11611 15668 11621
rect 15634 11543 15668 11549
rect 15634 11475 15668 11477
rect 15634 11439 15668 11441
rect 15634 11367 15668 11373
rect 15634 11295 15668 11305
rect 15634 11223 15668 11237
rect 15634 11151 15668 11169
rect 15634 11066 15668 11101
rect 15722 13039 15756 13074
rect 15722 12971 15756 12989
rect 15722 12903 15756 12917
rect 15722 12835 15756 12845
rect 15722 12767 15756 12773
rect 15722 12699 15756 12701
rect 15722 12663 15756 12665
rect 15722 12591 15756 12597
rect 15722 12519 15756 12529
rect 15722 12447 15756 12461
rect 15722 12375 15756 12393
rect 15722 12303 15756 12325
rect 15722 12231 15756 12257
rect 15722 12159 15756 12189
rect 15722 12087 15756 12121
rect 15722 12019 15756 12053
rect 15722 11951 15756 11981
rect 15722 11883 15756 11909
rect 15722 11815 15756 11837
rect 15722 11747 15756 11765
rect 15722 11679 15756 11693
rect 15722 11611 15756 11621
rect 15722 11543 15756 11549
rect 15722 11475 15756 11477
rect 15722 11439 15756 11441
rect 15722 11367 15756 11373
rect 15722 11295 15756 11305
rect 15722 11223 15756 11237
rect 15722 11151 15756 11169
rect 15722 11066 15756 11101
rect 15810 13039 15844 13074
rect 15810 12971 15844 12989
rect 15810 12903 15844 12917
rect 15810 12835 15844 12845
rect 15810 12767 15844 12773
rect 15810 12699 15844 12701
rect 15810 12663 15844 12665
rect 15810 12591 15844 12597
rect 15810 12519 15844 12529
rect 15810 12447 15844 12461
rect 15810 12375 15844 12393
rect 15810 12303 15844 12325
rect 15810 12231 15844 12257
rect 15810 12159 15844 12189
rect 15810 12087 15844 12121
rect 15810 12019 15844 12053
rect 15810 11951 15844 11981
rect 15810 11883 15844 11909
rect 15810 11815 15844 11837
rect 15810 11747 15844 11765
rect 15810 11679 15844 11693
rect 15810 11611 15844 11621
rect 15810 11543 15844 11549
rect 15810 11475 15844 11477
rect 15810 11439 15844 11441
rect 15810 11367 15844 11373
rect 15810 11295 15844 11305
rect 15810 11223 15844 11237
rect 15810 11151 15844 11169
rect 15810 11066 15844 11101
rect 15898 13039 15932 13074
rect 15898 12971 15932 12989
rect 15898 12903 15932 12917
rect 15898 12835 15932 12845
rect 15898 12767 15932 12773
rect 15898 12699 15932 12701
rect 15898 12663 15932 12665
rect 15898 12591 15932 12597
rect 15898 12519 15932 12529
rect 15898 12447 15932 12461
rect 15898 12375 15932 12393
rect 15898 12303 15932 12325
rect 15898 12231 15932 12257
rect 15898 12159 15932 12189
rect 15898 12087 15932 12121
rect 15898 12019 15932 12053
rect 15898 11951 15932 11981
rect 15898 11883 15932 11909
rect 15898 11815 15932 11837
rect 15898 11747 15932 11765
rect 15898 11679 15932 11693
rect 15898 11611 15932 11621
rect 15898 11543 15932 11549
rect 15898 11475 15932 11477
rect 15898 11439 15932 11441
rect 15898 11367 15932 11373
rect 15898 11295 15932 11305
rect 15898 11223 15932 11237
rect 15898 11151 15932 11169
rect 15898 11066 15932 11101
rect 15986 13039 16020 13074
rect 15986 12971 16020 12989
rect 15986 12903 16020 12917
rect 15986 12835 16020 12845
rect 15986 12767 16020 12773
rect 15986 12699 16020 12701
rect 15986 12663 16020 12665
rect 15986 12591 16020 12597
rect 15986 12519 16020 12529
rect 15986 12447 16020 12461
rect 15986 12375 16020 12393
rect 15986 12303 16020 12325
rect 15986 12231 16020 12257
rect 15986 12159 16020 12189
rect 15986 12087 16020 12121
rect 15986 12019 16020 12053
rect 15986 11951 16020 11981
rect 15986 11883 16020 11909
rect 15986 11815 16020 11837
rect 15986 11747 16020 11765
rect 15986 11679 16020 11693
rect 15986 11611 16020 11621
rect 15986 11543 16020 11549
rect 15986 11475 16020 11477
rect 15986 11439 16020 11441
rect 15986 11367 16020 11373
rect 15986 11295 16020 11305
rect 15986 11223 16020 11237
rect 15986 11151 16020 11169
rect 15986 11066 16020 11101
rect 16074 13039 16108 13074
rect 16074 12971 16108 12989
rect 16074 12903 16108 12917
rect 16074 12835 16108 12845
rect 16074 12767 16108 12773
rect 16074 12699 16108 12701
rect 16074 12663 16108 12665
rect 16074 12591 16108 12597
rect 16074 12519 16108 12529
rect 16074 12447 16108 12461
rect 16074 12375 16108 12393
rect 16074 12303 16108 12325
rect 16074 12231 16108 12257
rect 16074 12159 16108 12189
rect 16074 12087 16108 12121
rect 16074 12019 16108 12053
rect 16074 11951 16108 11981
rect 16074 11883 16108 11909
rect 16074 11815 16108 11837
rect 16074 11747 16108 11765
rect 16074 11679 16108 11693
rect 16074 11611 16108 11621
rect 16074 11543 16108 11549
rect 16074 11475 16108 11477
rect 16074 11439 16108 11441
rect 16074 11367 16108 11373
rect 16074 11295 16108 11305
rect 16074 11223 16108 11237
rect 16074 11151 16108 11169
rect 16074 11066 16108 11101
rect 16162 13039 16196 13074
rect 16162 12971 16196 12989
rect 16162 12903 16196 12917
rect 16162 12835 16196 12845
rect 16162 12767 16196 12773
rect 16162 12699 16196 12701
rect 16162 12663 16196 12665
rect 16162 12591 16196 12597
rect 16162 12519 16196 12529
rect 16162 12447 16196 12461
rect 16162 12375 16196 12393
rect 16162 12303 16196 12325
rect 16162 12231 16196 12257
rect 16162 12159 16196 12189
rect 16162 12087 16196 12121
rect 16162 12019 16196 12053
rect 16162 11951 16196 11981
rect 16162 11883 16196 11909
rect 16162 11815 16196 11837
rect 16162 11747 16196 11765
rect 16162 11679 16196 11693
rect 16162 11611 16196 11621
rect 16162 11543 16196 11549
rect 16162 11475 16196 11477
rect 16162 11439 16196 11441
rect 16162 11367 16196 11373
rect 16162 11295 16196 11305
rect 16162 11223 16196 11237
rect 16162 11151 16196 11169
rect 16162 11066 16196 11101
rect 16250 13039 16284 13074
rect 16250 12971 16284 12989
rect 16250 12903 16284 12917
rect 16250 12835 16284 12845
rect 16250 12767 16284 12773
rect 16250 12699 16284 12701
rect 16250 12663 16284 12665
rect 16250 12591 16284 12597
rect 16250 12519 16284 12529
rect 16250 12447 16284 12461
rect 16250 12375 16284 12393
rect 16250 12303 16284 12325
rect 16250 12231 16284 12257
rect 16250 12159 16284 12189
rect 16250 12087 16284 12121
rect 16250 12019 16284 12053
rect 16250 11951 16284 11981
rect 16250 11883 16284 11909
rect 16250 11815 16284 11837
rect 16250 11747 16284 11765
rect 16250 11679 16284 11693
rect 16250 11611 16284 11621
rect 16250 11543 16284 11549
rect 16250 11475 16284 11477
rect 16250 11439 16284 11441
rect 16250 11367 16284 11373
rect 16250 11295 16284 11305
rect 16250 11223 16284 11237
rect 16250 11151 16284 11169
rect 16250 11066 16284 11101
rect 16338 13039 16372 13074
rect 16338 12971 16372 12989
rect 16338 12903 16372 12917
rect 16338 12835 16372 12845
rect 16338 12767 16372 12773
rect 16338 12699 16372 12701
rect 16338 12663 16372 12665
rect 16338 12591 16372 12597
rect 16338 12519 16372 12529
rect 16338 12447 16372 12461
rect 16338 12375 16372 12393
rect 16338 12303 16372 12325
rect 16338 12231 16372 12257
rect 16338 12159 16372 12189
rect 16338 12087 16372 12121
rect 16338 12019 16372 12053
rect 16338 11951 16372 11981
rect 16338 11883 16372 11909
rect 16338 11815 16372 11837
rect 16338 11747 16372 11765
rect 16338 11679 16372 11693
rect 16338 11611 16372 11621
rect 16338 11543 16372 11549
rect 16338 11475 16372 11477
rect 16338 11439 16372 11441
rect 16338 11367 16372 11373
rect 16338 11295 16372 11305
rect 16338 11223 16372 11237
rect 16338 11151 16372 11169
rect 16338 11066 16372 11101
rect 16426 13039 16460 13074
rect 16426 12971 16460 12989
rect 16426 12903 16460 12917
rect 16426 12835 16460 12845
rect 16426 12767 16460 12773
rect 16426 12699 16460 12701
rect 16426 12663 16460 12665
rect 16426 12591 16460 12597
rect 16426 12519 16460 12529
rect 16426 12447 16460 12461
rect 16426 12375 16460 12393
rect 16426 12303 16460 12325
rect 16426 12231 16460 12257
rect 16426 12159 16460 12189
rect 16426 12087 16460 12121
rect 16426 12019 16460 12053
rect 16426 11951 16460 11981
rect 16426 11883 16460 11909
rect 16426 11815 16460 11837
rect 16426 11747 16460 11765
rect 16426 11679 16460 11693
rect 16426 11611 16460 11621
rect 16426 11543 16460 11549
rect 16426 11475 16460 11477
rect 16426 11439 16460 11441
rect 16426 11367 16460 11373
rect 16426 11295 16460 11305
rect 16426 11223 16460 11237
rect 16426 11151 16460 11169
rect 16426 11066 16460 11101
rect 16514 13039 16548 13074
rect 16514 12971 16548 12989
rect 16514 12903 16548 12917
rect 16514 12835 16548 12845
rect 16514 12767 16548 12773
rect 16514 12699 16548 12701
rect 16514 12663 16548 12665
rect 16514 12591 16548 12597
rect 16514 12519 16548 12529
rect 16514 12447 16548 12461
rect 16514 12375 16548 12393
rect 16514 12303 16548 12325
rect 16514 12231 16548 12257
rect 16514 12159 16548 12189
rect 16514 12087 16548 12121
rect 16514 12019 16548 12053
rect 16514 11951 16548 11981
rect 16514 11883 16548 11909
rect 16514 11815 16548 11837
rect 16514 11747 16548 11765
rect 16514 11679 16548 11693
rect 16514 11611 16548 11621
rect 16514 11543 16548 11549
rect 16514 11475 16548 11477
rect 16514 11439 16548 11441
rect 16514 11367 16548 11373
rect 16514 11295 16548 11305
rect 16514 11223 16548 11237
rect 16514 11151 16548 11169
rect 16514 11066 16548 11101
rect 16602 13039 16636 13074
rect 16602 12971 16636 12989
rect 16602 12903 16636 12917
rect 16602 12835 16636 12845
rect 16602 12767 16636 12773
rect 16602 12699 16636 12701
rect 16602 12663 16636 12665
rect 16602 12591 16636 12597
rect 16602 12519 16636 12529
rect 16602 12447 16636 12461
rect 16602 12375 16636 12393
rect 16602 12303 16636 12325
rect 16602 12231 16636 12257
rect 16602 12159 16636 12189
rect 16602 12087 16636 12121
rect 16602 12019 16636 12053
rect 16602 11951 16636 11981
rect 16602 11883 16636 11909
rect 16602 11815 16636 11837
rect 16602 11747 16636 11765
rect 16602 11679 16636 11693
rect 16602 11611 16636 11621
rect 16602 11543 16636 11549
rect 16602 11475 16636 11477
rect 16602 11439 16636 11441
rect 16602 11367 16636 11373
rect 16602 11295 16636 11305
rect 16602 11223 16636 11237
rect 16602 11151 16636 11169
rect 16602 11066 16636 11101
rect 16690 13039 16724 13074
rect 16690 12971 16724 12989
rect 16690 12903 16724 12917
rect 16690 12835 16724 12845
rect 16690 12767 16724 12773
rect 16690 12699 16724 12701
rect 16690 12663 16724 12665
rect 16690 12591 16724 12597
rect 16690 12519 16724 12529
rect 16690 12447 16724 12461
rect 16690 12375 16724 12393
rect 16690 12303 16724 12325
rect 16690 12231 16724 12257
rect 16690 12159 16724 12189
rect 16690 12087 16724 12121
rect 16690 12019 16724 12053
rect 16690 11951 16724 11981
rect 16690 11883 16724 11909
rect 16690 11815 16724 11837
rect 16690 11747 16724 11765
rect 16690 11679 16724 11693
rect 16690 11611 16724 11621
rect 16690 11543 16724 11549
rect 16690 11475 16724 11477
rect 16690 11439 16724 11441
rect 16690 11367 16724 11373
rect 16690 11295 16724 11305
rect 16690 11223 16724 11237
rect 16690 11151 16724 11169
rect 16690 11066 16724 11101
rect 16778 13039 16812 13074
rect 16778 12971 16812 12989
rect 16778 12903 16812 12917
rect 16778 12835 16812 12845
rect 16778 12767 16812 12773
rect 16778 12699 16812 12701
rect 16778 12663 16812 12665
rect 16778 12591 16812 12597
rect 16778 12519 16812 12529
rect 16778 12447 16812 12461
rect 16778 12375 16812 12393
rect 16778 12303 16812 12325
rect 16778 12231 16812 12257
rect 16778 12159 16812 12189
rect 16778 12087 16812 12121
rect 16778 12019 16812 12053
rect 16778 11951 16812 11981
rect 16778 11883 16812 11909
rect 16778 11815 16812 11837
rect 16778 11747 16812 11765
rect 16778 11679 16812 11693
rect 16778 11611 16812 11621
rect 16778 11543 16812 11549
rect 16778 11475 16812 11477
rect 16778 11439 16812 11441
rect 16778 11367 16812 11373
rect 16778 11295 16812 11305
rect 16778 11223 16812 11237
rect 16778 11151 16812 11169
rect 16778 11066 16812 11101
rect 16866 13039 16900 13074
rect 16866 12971 16900 12989
rect 16866 12903 16900 12917
rect 16866 12835 16900 12845
rect 16866 12767 16900 12773
rect 16866 12699 16900 12701
rect 16866 12663 16900 12665
rect 16866 12591 16900 12597
rect 16866 12519 16900 12529
rect 16866 12447 16900 12461
rect 16866 12375 16900 12393
rect 16866 12303 16900 12325
rect 16866 12231 16900 12257
rect 16866 12159 16900 12189
rect 16866 12087 16900 12121
rect 16866 12019 16900 12053
rect 16866 11951 16900 11981
rect 16866 11883 16900 11909
rect 16866 11815 16900 11837
rect 16866 11747 16900 11765
rect 16866 11679 16900 11693
rect 16866 11611 16900 11621
rect 16866 11543 16900 11549
rect 16866 11475 16900 11477
rect 16866 11439 16900 11441
rect 16866 11367 16900 11373
rect 16866 11295 16900 11305
rect 16866 11223 16900 11237
rect 16866 11151 16900 11169
rect 16866 11066 16900 11101
rect 16954 13039 16988 13074
rect 16954 12971 16988 12989
rect 16954 12903 16988 12917
rect 16954 12835 16988 12845
rect 16954 12767 16988 12773
rect 16954 12699 16988 12701
rect 16954 12663 16988 12665
rect 16954 12591 16988 12597
rect 16954 12519 16988 12529
rect 16954 12447 16988 12461
rect 16954 12375 16988 12393
rect 16954 12303 16988 12325
rect 16954 12231 16988 12257
rect 16954 12159 16988 12189
rect 16954 12087 16988 12121
rect 16954 12019 16988 12053
rect 16954 11951 16988 11981
rect 16954 11883 16988 11909
rect 16954 11815 16988 11837
rect 16954 11747 16988 11765
rect 16954 11679 16988 11693
rect 16954 11611 16988 11621
rect 16954 11543 16988 11549
rect 16954 11475 16988 11477
rect 16954 11439 16988 11441
rect 16954 11367 16988 11373
rect 16954 11295 16988 11305
rect 16954 11223 16988 11237
rect 16954 11151 16988 11169
rect 16954 11066 16988 11101
rect 17042 13039 17076 13074
rect 17042 12971 17076 12989
rect 17042 12903 17076 12917
rect 17042 12835 17076 12845
rect 17042 12767 17076 12773
rect 17042 12699 17076 12701
rect 17042 12663 17076 12665
rect 17042 12591 17076 12597
rect 17042 12519 17076 12529
rect 17042 12447 17076 12461
rect 17042 12375 17076 12393
rect 17042 12303 17076 12325
rect 17042 12231 17076 12257
rect 17042 12159 17076 12189
rect 17042 12087 17076 12121
rect 17042 12019 17076 12053
rect 17042 11951 17076 11981
rect 17042 11883 17076 11909
rect 17042 11815 17076 11837
rect 17042 11747 17076 11765
rect 17042 11679 17076 11693
rect 17042 11611 17076 11621
rect 17042 11543 17076 11549
rect 17042 11475 17076 11477
rect 17042 11439 17076 11441
rect 17042 11367 17076 11373
rect 17042 11295 17076 11305
rect 17042 11223 17076 11237
rect 17042 11151 17076 11169
rect 17042 11066 17076 11101
rect 17130 13039 17164 13074
rect 17130 12971 17164 12989
rect 17130 12903 17164 12917
rect 17130 12835 17164 12845
rect 17130 12767 17164 12773
rect 17130 12699 17164 12701
rect 17130 12663 17164 12665
rect 17130 12591 17164 12597
rect 17130 12519 17164 12529
rect 17130 12447 17164 12461
rect 17130 12375 17164 12393
rect 17130 12303 17164 12325
rect 17130 12231 17164 12257
rect 17130 12159 17164 12189
rect 17130 12087 17164 12121
rect 17130 12019 17164 12053
rect 17130 11951 17164 11981
rect 17130 11883 17164 11909
rect 17130 11815 17164 11837
rect 17130 11747 17164 11765
rect 17130 11679 17164 11693
rect 17130 11611 17164 11621
rect 17130 11543 17164 11549
rect 17130 11475 17164 11477
rect 17130 11439 17164 11441
rect 17130 11367 17164 11373
rect 17130 11295 17164 11305
rect 17130 11223 17164 11237
rect 17130 11151 17164 11169
rect 17130 11066 17164 11101
rect 17218 13039 17252 13074
rect 17218 12971 17252 12989
rect 17218 12903 17252 12917
rect 17218 12835 17252 12845
rect 17218 12767 17252 12773
rect 17218 12699 17252 12701
rect 17218 12663 17252 12665
rect 17218 12591 17252 12597
rect 17218 12519 17252 12529
rect 17218 12447 17252 12461
rect 17218 12375 17252 12393
rect 17218 12303 17252 12325
rect 17218 12231 17252 12257
rect 17218 12159 17252 12189
rect 17218 12087 17252 12121
rect 17218 12019 17252 12053
rect 17218 11951 17252 11981
rect 17218 11883 17252 11909
rect 17218 11815 17252 11837
rect 17218 11747 17252 11765
rect 17218 11679 17252 11693
rect 17218 11611 17252 11621
rect 17218 11543 17252 11549
rect 17218 11475 17252 11477
rect 17218 11439 17252 11441
rect 17218 11367 17252 11373
rect 17218 11295 17252 11305
rect 17218 11223 17252 11237
rect 17218 11151 17252 11169
rect 17218 11066 17252 11101
rect 17306 13039 17340 13074
rect 17306 12971 17340 12989
rect 17306 12903 17340 12917
rect 17306 12835 17340 12845
rect 17306 12767 17340 12773
rect 17306 12699 17340 12701
rect 17306 12663 17340 12665
rect 17306 12591 17340 12597
rect 17306 12519 17340 12529
rect 17306 12447 17340 12461
rect 17306 12375 17340 12393
rect 17306 12303 17340 12325
rect 17306 12231 17340 12257
rect 17306 12159 17340 12189
rect 17306 12087 17340 12121
rect 17306 12019 17340 12053
rect 17306 11951 17340 11981
rect 17306 11883 17340 11909
rect 17306 11815 17340 11837
rect 17306 11747 17340 11765
rect 17306 11679 17340 11693
rect 17306 11611 17340 11621
rect 17306 11543 17340 11549
rect 17306 11475 17340 11477
rect 17306 11439 17340 11441
rect 17306 11367 17340 11373
rect 17306 11295 17340 11305
rect 17306 11223 17340 11237
rect 17306 11151 17340 11169
rect 17306 11066 17340 11101
rect 17394 13039 17428 13074
rect 17394 12971 17428 12989
rect 17394 12903 17428 12917
rect 17394 12835 17428 12845
rect 17394 12767 17428 12773
rect 17394 12699 17428 12701
rect 17394 12663 17428 12665
rect 17394 12591 17428 12597
rect 17394 12519 17428 12529
rect 17394 12447 17428 12461
rect 17394 12375 17428 12393
rect 17394 12303 17428 12325
rect 17394 12231 17428 12257
rect 17394 12159 17428 12189
rect 17394 12087 17428 12121
rect 17394 12019 17428 12053
rect 17394 11951 17428 11981
rect 17394 11883 17428 11909
rect 17394 11815 17428 11837
rect 17394 11747 17428 11765
rect 17394 11679 17428 11693
rect 17394 11611 17428 11621
rect 17394 11543 17428 11549
rect 17394 11475 17428 11477
rect 17394 11439 17428 11441
rect 17394 11367 17428 11373
rect 17394 11295 17428 11305
rect 17394 11223 17428 11237
rect 17394 11151 17428 11169
rect 17394 11066 17428 11101
rect 17482 13039 17516 13074
rect 17482 12971 17516 12989
rect 17482 12903 17516 12917
rect 17482 12835 17516 12845
rect 17482 12767 17516 12773
rect 17482 12699 17516 12701
rect 17482 12663 17516 12665
rect 17482 12591 17516 12597
rect 17482 12519 17516 12529
rect 17482 12447 17516 12461
rect 17482 12375 17516 12393
rect 17482 12303 17516 12325
rect 17482 12231 17516 12257
rect 17482 12159 17516 12189
rect 17482 12087 17516 12121
rect 17482 12019 17516 12053
rect 17482 11951 17516 11981
rect 17482 11883 17516 11909
rect 17482 11815 17516 11837
rect 17482 11747 17516 11765
rect 17482 11679 17516 11693
rect 17482 11611 17516 11621
rect 17482 11543 17516 11549
rect 17482 11475 17516 11477
rect 17482 11439 17516 11441
rect 17482 11367 17516 11373
rect 17482 11295 17516 11305
rect 17482 11223 17516 11237
rect 17482 11151 17516 11169
rect 17482 11066 17516 11101
rect 17728 13051 17785 13085
rect 17819 13051 17870 13085
rect 17728 13017 17870 13051
rect 17728 12983 17785 13017
rect 17819 12983 17870 13017
rect 17728 12949 17870 12983
rect 17728 12915 17785 12949
rect 17819 12915 17870 12949
rect 17728 12881 17870 12915
rect 17728 12847 17785 12881
rect 17819 12847 17870 12881
rect 17728 12813 17870 12847
rect 17728 12779 17785 12813
rect 17819 12779 17870 12813
rect 17728 12745 17870 12779
rect 17728 12711 17785 12745
rect 17819 12711 17870 12745
rect 17728 12677 17870 12711
rect 17728 12643 17785 12677
rect 17819 12643 17870 12677
rect 17728 12609 17870 12643
rect 17728 12575 17785 12609
rect 17819 12575 17870 12609
rect 17728 12541 17870 12575
rect 17728 12507 17785 12541
rect 17819 12507 17870 12541
rect 17728 12473 17870 12507
rect 17728 12439 17785 12473
rect 17819 12439 17870 12473
rect 17728 12405 17870 12439
rect 17728 12371 17785 12405
rect 17819 12371 17870 12405
rect 17728 12337 17870 12371
rect 17728 12303 17785 12337
rect 17819 12303 17870 12337
rect 17728 12269 17870 12303
rect 17728 12235 17785 12269
rect 17819 12235 17870 12269
rect 17728 12201 17870 12235
rect 17728 12167 17785 12201
rect 17819 12167 17870 12201
rect 17728 12133 17870 12167
rect 17728 12099 17785 12133
rect 17819 12099 17870 12133
rect 17728 12065 17870 12099
rect 17728 12031 17785 12065
rect 17819 12031 17870 12065
rect 17728 11997 17870 12031
rect 17728 11963 17785 11997
rect 17819 11963 17870 11997
rect 17728 11929 17870 11963
rect 17728 11895 17785 11929
rect 17819 11895 17870 11929
rect 17728 11861 17870 11895
rect 17728 11827 17785 11861
rect 17819 11827 17870 11861
rect 17728 11793 17870 11827
rect 17728 11759 17785 11793
rect 17819 11759 17870 11793
rect 17728 11725 17870 11759
rect 17728 11691 17785 11725
rect 17819 11691 17870 11725
rect 17728 11657 17870 11691
rect 17728 11623 17785 11657
rect 17819 11623 17870 11657
rect 17728 11589 17870 11623
rect 17728 11555 17785 11589
rect 17819 11555 17870 11589
rect 17728 11521 17870 11555
rect 17728 11487 17785 11521
rect 17819 11487 17870 11521
rect 17728 11453 17870 11487
rect 17728 11419 17785 11453
rect 17819 11419 17870 11453
rect 17728 11385 17870 11419
rect 17728 11351 17785 11385
rect 17819 11351 17870 11385
rect 17728 11317 17870 11351
rect 17728 11283 17785 11317
rect 17819 11283 17870 11317
rect 17728 11249 17870 11283
rect 17728 11215 17785 11249
rect 17819 11215 17870 11249
rect 17728 11181 17870 11215
rect 17728 11147 17785 11181
rect 17819 11147 17870 11181
rect 17728 11113 17870 11147
rect 17728 11079 17785 11113
rect 17819 11079 17870 11113
rect 13074 11002 13122 11036
rect 13156 11002 13209 11036
rect 17728 11045 17870 11079
rect 13074 10968 13209 11002
rect 13497 11000 13572 11020
rect 13847 11000 13922 11014
rect 14205 11000 14280 11017
rect 14553 11000 14628 11017
rect 14904 11000 14979 11017
rect 15255 11000 15330 11016
rect 15606 11000 15681 11014
rect 15961 11000 16036 11017
rect 16311 11000 16386 11013
rect 16665 11000 16740 11015
rect 17015 11000 17090 11013
rect 13074 10934 13122 10968
rect 13156 10934 13209 10968
rect 13074 10900 13209 10934
rect 13074 10866 13122 10900
rect 13156 10866 13209 10900
rect 13074 10832 13209 10866
rect 13074 10798 13122 10832
rect 13156 10798 13209 10832
rect 13467 10996 17158 11000
rect 13467 10962 13517 10996
rect 13551 10993 17158 10996
rect 13551 10990 14225 10993
rect 13551 10962 13867 10990
rect 13467 10956 13867 10962
rect 13901 10959 14225 10990
rect 14259 10959 14573 10993
rect 14607 10959 14924 10993
rect 14958 10992 15981 10993
rect 14958 10959 15275 10992
rect 13901 10958 15275 10959
rect 15309 10990 15981 10992
rect 15309 10958 15626 10990
rect 13901 10956 15626 10958
rect 15660 10959 15981 10990
rect 16015 10991 17158 10993
rect 16015 10989 16685 10991
rect 16015 10959 16331 10989
rect 15660 10956 16331 10959
rect 13467 10955 16331 10956
rect 16365 10957 16685 10989
rect 16719 10989 17158 10991
rect 16719 10957 17035 10989
rect 16365 10955 17035 10957
rect 17069 10955 17158 10989
rect 13467 10931 17158 10955
rect 17352 10971 17472 11024
rect 17352 10937 17395 10971
rect 17429 10937 17472 10971
rect 13467 10861 13597 10931
rect 17352 10894 17472 10937
rect 17728 11011 17785 11045
rect 17819 11011 17870 11045
rect 17728 10977 17870 11011
rect 17728 10943 17785 10977
rect 17819 10943 17870 10977
rect 17728 10909 17870 10943
rect 13467 10827 13514 10861
rect 13548 10827 13597 10861
rect 13467 10804 13597 10827
rect 17342 10846 17482 10894
rect 17342 10812 17395 10846
rect 17429 10812 17482 10846
rect 13074 10738 13209 10798
rect 17342 10774 17482 10812
rect 17728 10875 17785 10909
rect 17819 10875 17870 10909
rect 17728 10841 17870 10875
rect 17728 10807 17785 10841
rect 17819 10807 17870 10841
rect 17728 10738 17870 10807
rect 13074 10701 17870 10738
rect 13074 10693 14503 10701
rect 14537 10693 14575 10701
rect 14609 10693 14647 10701
rect 14681 10693 17870 10701
rect 13074 10659 13371 10693
rect 13405 10659 13439 10693
rect 13473 10659 13507 10693
rect 13541 10659 13575 10693
rect 13609 10659 13643 10693
rect 13677 10659 13711 10693
rect 13745 10659 13779 10693
rect 13813 10659 13847 10693
rect 13881 10659 13915 10693
rect 13949 10659 13983 10693
rect 14017 10659 14051 10693
rect 14085 10659 14119 10693
rect 14153 10659 14187 10693
rect 14221 10659 14255 10693
rect 14289 10659 14323 10693
rect 14357 10659 14391 10693
rect 14425 10659 14459 10693
rect 14493 10667 14503 10693
rect 14561 10667 14575 10693
rect 14629 10667 14647 10693
rect 14493 10659 14527 10667
rect 14561 10659 14595 10667
rect 14629 10659 14663 10667
rect 14697 10659 14731 10693
rect 14765 10659 14799 10693
rect 14833 10659 14867 10693
rect 14901 10659 14935 10693
rect 14969 10659 15003 10693
rect 15037 10659 15071 10693
rect 15105 10659 15139 10693
rect 15173 10659 15207 10693
rect 15241 10659 15275 10693
rect 15309 10659 15343 10693
rect 15377 10659 15411 10693
rect 15445 10659 15479 10693
rect 15513 10659 15547 10693
rect 15581 10659 15615 10693
rect 15649 10659 15683 10693
rect 15717 10659 15751 10693
rect 15785 10659 15819 10693
rect 15853 10659 15887 10693
rect 15921 10659 15955 10693
rect 15989 10659 16023 10693
rect 16057 10659 16091 10693
rect 16125 10659 16159 10693
rect 16193 10659 16227 10693
rect 16261 10659 16295 10693
rect 16329 10659 16363 10693
rect 16397 10659 16431 10693
rect 16465 10659 16499 10693
rect 16533 10659 16567 10693
rect 16601 10659 16635 10693
rect 16669 10659 16703 10693
rect 16737 10659 16771 10693
rect 16805 10659 16839 10693
rect 16873 10659 16907 10693
rect 16941 10659 16975 10693
rect 17009 10659 17043 10693
rect 17077 10659 17111 10693
rect 17145 10659 17179 10693
rect 17213 10659 17247 10693
rect 17281 10659 17315 10693
rect 17349 10659 17383 10693
rect 17417 10659 17451 10693
rect 17485 10659 17519 10693
rect 17553 10659 17587 10693
rect 17621 10659 17870 10693
rect 13074 10610 17870 10659
rect 13861 10532 17005 10610
rect 13850 9654 17008 10532
rect 13850 8972 13929 9654
rect 16915 8972 17008 9654
rect 13850 8882 17008 8972
<< viali >>
rect 14128 27701 16394 28815
rect 13065 24564 13099 24598
rect 13137 24564 13171 24598
rect 13209 24564 13243 24598
rect 13281 24564 13315 24598
rect 13353 24564 13387 24598
rect 13425 24564 13459 24598
rect 16496 24564 16530 24598
rect 16568 24564 16602 24598
rect 16640 24564 16674 24598
rect 16712 24564 16746 24598
rect 16784 24564 16818 24598
rect 16856 24564 16890 24598
rect 16806 24078 16840 24112
rect 16998 24078 17032 24112
rect 17190 24078 17224 24112
rect 17382 24078 17416 24112
rect 17574 24078 17608 24112
rect 13095 23884 13129 23918
rect 13167 23884 13201 23918
rect 13239 23884 13273 23918
rect 13311 23884 13345 23918
rect 13383 23884 13417 23918
rect 13455 23884 13489 23918
rect 14326 23884 14360 23918
rect 14398 23884 14432 23918
rect 14470 23884 14504 23918
rect 14542 23884 14576 23918
rect 14614 23884 14648 23918
rect 14686 23884 14720 23918
rect 13111 23417 13289 23523
rect 16307 23442 16413 23548
rect 14114 23188 14148 23222
rect 14306 23188 14340 23222
rect 14498 23188 14532 23222
rect 14690 23188 14724 23222
rect 13504 22016 13538 22050
rect 13504 21944 13538 21978
rect 13504 21872 13538 21906
rect 13504 21800 13538 21834
rect 13504 21728 13538 21762
rect 13504 21656 13538 21690
rect 13504 21485 13538 21519
rect 13504 21413 13538 21447
rect 13504 21341 13538 21375
rect 13504 21269 13538 21303
rect 13504 21197 13538 21231
rect 13504 21125 13538 21159
rect 13970 23085 14004 23103
rect 13970 23069 14004 23085
rect 13970 23017 14004 23031
rect 13970 22997 14004 23017
rect 13970 22949 14004 22959
rect 13970 22925 14004 22949
rect 13970 22881 14004 22887
rect 13970 22853 14004 22881
rect 13970 22813 14004 22815
rect 13970 22781 14004 22813
rect 13970 22711 14004 22743
rect 13970 22709 14004 22711
rect 13970 22643 14004 22671
rect 13970 22637 14004 22643
rect 13970 22575 14004 22599
rect 13970 22565 14004 22575
rect 13970 22507 14004 22527
rect 13970 22493 14004 22507
rect 13970 22439 14004 22455
rect 13970 22421 14004 22439
rect 13970 22371 14004 22383
rect 13970 22349 14004 22371
rect 13970 22303 14004 22311
rect 13970 22277 14004 22303
rect 13970 22235 14004 22239
rect 13970 22205 14004 22235
rect 13970 22133 14004 22167
rect 13970 22065 14004 22095
rect 13970 22061 14004 22065
rect 13970 21997 14004 22023
rect 13970 21989 14004 21997
rect 13970 21929 14004 21951
rect 13970 21917 14004 21929
rect 13970 21861 14004 21879
rect 13970 21845 14004 21861
rect 13970 21793 14004 21807
rect 13970 21773 14004 21793
rect 13970 21725 14004 21735
rect 13970 21701 14004 21725
rect 13970 21657 14004 21663
rect 13970 21629 14004 21657
rect 13970 21589 14004 21591
rect 13970 21557 14004 21589
rect 13970 21487 14004 21519
rect 13970 21485 14004 21487
rect 13970 21419 14004 21447
rect 13970 21413 14004 21419
rect 13970 21351 14004 21375
rect 13970 21341 14004 21351
rect 13970 21283 14004 21303
rect 13970 21269 14004 21283
rect 13970 21215 14004 21231
rect 13970 21197 14004 21215
rect 14066 23085 14100 23103
rect 14066 23069 14100 23085
rect 14066 23017 14100 23031
rect 14066 22997 14100 23017
rect 14066 22949 14100 22959
rect 14066 22925 14100 22949
rect 14066 22881 14100 22887
rect 14066 22853 14100 22881
rect 14066 22813 14100 22815
rect 14066 22781 14100 22813
rect 14066 22711 14100 22743
rect 14066 22709 14100 22711
rect 14066 22643 14100 22671
rect 14066 22637 14100 22643
rect 14066 22575 14100 22599
rect 14066 22565 14100 22575
rect 14066 22507 14100 22527
rect 14066 22493 14100 22507
rect 14066 22439 14100 22455
rect 14066 22421 14100 22439
rect 14066 22371 14100 22383
rect 14066 22349 14100 22371
rect 14066 22303 14100 22311
rect 14066 22277 14100 22303
rect 14066 22235 14100 22239
rect 14066 22205 14100 22235
rect 14066 22133 14100 22167
rect 14066 22065 14100 22095
rect 14066 22061 14100 22065
rect 14066 21997 14100 22023
rect 14066 21989 14100 21997
rect 14066 21929 14100 21951
rect 14066 21917 14100 21929
rect 14066 21861 14100 21879
rect 14066 21845 14100 21861
rect 14066 21793 14100 21807
rect 14066 21773 14100 21793
rect 14066 21725 14100 21735
rect 14066 21701 14100 21725
rect 14066 21657 14100 21663
rect 14066 21629 14100 21657
rect 14066 21589 14100 21591
rect 14066 21557 14100 21589
rect 14066 21487 14100 21519
rect 14066 21485 14100 21487
rect 14066 21419 14100 21447
rect 14066 21413 14100 21419
rect 14066 21351 14100 21375
rect 14066 21341 14100 21351
rect 14066 21283 14100 21303
rect 14066 21269 14100 21283
rect 14066 21215 14100 21231
rect 14066 21197 14100 21215
rect 14162 23085 14196 23103
rect 14162 23069 14196 23085
rect 14162 23017 14196 23031
rect 14162 22997 14196 23017
rect 14162 22949 14196 22959
rect 14162 22925 14196 22949
rect 14162 22881 14196 22887
rect 14162 22853 14196 22881
rect 14162 22813 14196 22815
rect 14162 22781 14196 22813
rect 14162 22711 14196 22743
rect 14162 22709 14196 22711
rect 14162 22643 14196 22671
rect 14162 22637 14196 22643
rect 14162 22575 14196 22599
rect 14162 22565 14196 22575
rect 14162 22507 14196 22527
rect 14162 22493 14196 22507
rect 14162 22439 14196 22455
rect 14162 22421 14196 22439
rect 14162 22371 14196 22383
rect 14162 22349 14196 22371
rect 14162 22303 14196 22311
rect 14162 22277 14196 22303
rect 14162 22235 14196 22239
rect 14162 22205 14196 22235
rect 14162 22133 14196 22167
rect 14162 22065 14196 22095
rect 14162 22061 14196 22065
rect 14162 21997 14196 22023
rect 14162 21989 14196 21997
rect 14162 21929 14196 21951
rect 14162 21917 14196 21929
rect 14162 21861 14196 21879
rect 14162 21845 14196 21861
rect 14162 21793 14196 21807
rect 14162 21773 14196 21793
rect 14162 21725 14196 21735
rect 14162 21701 14196 21725
rect 14162 21657 14196 21663
rect 14162 21629 14196 21657
rect 14162 21589 14196 21591
rect 14162 21557 14196 21589
rect 14162 21487 14196 21519
rect 14162 21485 14196 21487
rect 14162 21419 14196 21447
rect 14162 21413 14196 21419
rect 14162 21351 14196 21375
rect 14162 21341 14196 21351
rect 14162 21283 14196 21303
rect 14162 21269 14196 21283
rect 14162 21215 14196 21231
rect 14162 21197 14196 21215
rect 14258 23085 14292 23103
rect 14258 23069 14292 23085
rect 14258 23017 14292 23031
rect 14258 22997 14292 23017
rect 14258 22949 14292 22959
rect 14258 22925 14292 22949
rect 14258 22881 14292 22887
rect 14258 22853 14292 22881
rect 14258 22813 14292 22815
rect 14258 22781 14292 22813
rect 14258 22711 14292 22743
rect 14258 22709 14292 22711
rect 14258 22643 14292 22671
rect 14258 22637 14292 22643
rect 14258 22575 14292 22599
rect 14258 22565 14292 22575
rect 14258 22507 14292 22527
rect 14258 22493 14292 22507
rect 14258 22439 14292 22455
rect 14258 22421 14292 22439
rect 14258 22371 14292 22383
rect 14258 22349 14292 22371
rect 14258 22303 14292 22311
rect 14258 22277 14292 22303
rect 14258 22235 14292 22239
rect 14258 22205 14292 22235
rect 14258 22133 14292 22167
rect 14258 22065 14292 22095
rect 14258 22061 14292 22065
rect 14258 21997 14292 22023
rect 14258 21989 14292 21997
rect 14258 21929 14292 21951
rect 14258 21917 14292 21929
rect 14258 21861 14292 21879
rect 14258 21845 14292 21861
rect 14258 21793 14292 21807
rect 14258 21773 14292 21793
rect 14258 21725 14292 21735
rect 14258 21701 14292 21725
rect 14258 21657 14292 21663
rect 14258 21629 14292 21657
rect 14258 21589 14292 21591
rect 14258 21557 14292 21589
rect 14258 21487 14292 21519
rect 14258 21485 14292 21487
rect 14258 21419 14292 21447
rect 14258 21413 14292 21419
rect 14258 21351 14292 21375
rect 14258 21341 14292 21351
rect 14258 21283 14292 21303
rect 14258 21269 14292 21283
rect 14258 21215 14292 21231
rect 14258 21197 14292 21215
rect 14354 23085 14388 23103
rect 14354 23069 14388 23085
rect 14354 23017 14388 23031
rect 14354 22997 14388 23017
rect 14354 22949 14388 22959
rect 14354 22925 14388 22949
rect 14354 22881 14388 22887
rect 14354 22853 14388 22881
rect 14354 22813 14388 22815
rect 14354 22781 14388 22813
rect 14354 22711 14388 22743
rect 14354 22709 14388 22711
rect 14354 22643 14388 22671
rect 14354 22637 14388 22643
rect 14354 22575 14388 22599
rect 14354 22565 14388 22575
rect 14354 22507 14388 22527
rect 14354 22493 14388 22507
rect 14354 22439 14388 22455
rect 14354 22421 14388 22439
rect 14354 22371 14388 22383
rect 14354 22349 14388 22371
rect 14354 22303 14388 22311
rect 14354 22277 14388 22303
rect 14354 22235 14388 22239
rect 14354 22205 14388 22235
rect 14354 22133 14388 22167
rect 14354 22065 14388 22095
rect 14354 22061 14388 22065
rect 14354 21997 14388 22023
rect 14354 21989 14388 21997
rect 14354 21929 14388 21951
rect 14354 21917 14388 21929
rect 14354 21861 14388 21879
rect 14354 21845 14388 21861
rect 14354 21793 14388 21807
rect 14354 21773 14388 21793
rect 14354 21725 14388 21735
rect 14354 21701 14388 21725
rect 14354 21657 14388 21663
rect 14354 21629 14388 21657
rect 14354 21589 14388 21591
rect 14354 21557 14388 21589
rect 14354 21487 14388 21519
rect 14354 21485 14388 21487
rect 14354 21419 14388 21447
rect 14354 21413 14388 21419
rect 14354 21351 14388 21375
rect 14354 21341 14388 21351
rect 14354 21283 14388 21303
rect 14354 21269 14388 21283
rect 14354 21215 14388 21231
rect 14354 21197 14388 21215
rect 14450 23085 14484 23103
rect 14450 23069 14484 23085
rect 14450 23017 14484 23031
rect 14450 22997 14484 23017
rect 14450 22949 14484 22959
rect 14450 22925 14484 22949
rect 14450 22881 14484 22887
rect 14450 22853 14484 22881
rect 14450 22813 14484 22815
rect 14450 22781 14484 22813
rect 14450 22711 14484 22743
rect 14450 22709 14484 22711
rect 14450 22643 14484 22671
rect 14450 22637 14484 22643
rect 14450 22575 14484 22599
rect 14450 22565 14484 22575
rect 14450 22507 14484 22527
rect 14450 22493 14484 22507
rect 14450 22439 14484 22455
rect 14450 22421 14484 22439
rect 14450 22371 14484 22383
rect 14450 22349 14484 22371
rect 14450 22303 14484 22311
rect 14450 22277 14484 22303
rect 14450 22235 14484 22239
rect 14450 22205 14484 22235
rect 14450 22133 14484 22167
rect 14450 22065 14484 22095
rect 14450 22061 14484 22065
rect 14450 21997 14484 22023
rect 14450 21989 14484 21997
rect 14450 21929 14484 21951
rect 14450 21917 14484 21929
rect 14450 21861 14484 21879
rect 14450 21845 14484 21861
rect 14450 21793 14484 21807
rect 14450 21773 14484 21793
rect 14450 21725 14484 21735
rect 14450 21701 14484 21725
rect 14450 21657 14484 21663
rect 14450 21629 14484 21657
rect 14450 21589 14484 21591
rect 14450 21557 14484 21589
rect 14450 21487 14484 21519
rect 14450 21485 14484 21487
rect 14450 21419 14484 21447
rect 14450 21413 14484 21419
rect 14450 21351 14484 21375
rect 14450 21341 14484 21351
rect 14450 21283 14484 21303
rect 14450 21269 14484 21283
rect 14450 21215 14484 21231
rect 14450 21197 14484 21215
rect 14546 23085 14580 23103
rect 14546 23069 14580 23085
rect 14546 23017 14580 23031
rect 14546 22997 14580 23017
rect 14546 22949 14580 22959
rect 14546 22925 14580 22949
rect 14546 22881 14580 22887
rect 14546 22853 14580 22881
rect 14546 22813 14580 22815
rect 14546 22781 14580 22813
rect 14546 22711 14580 22743
rect 14546 22709 14580 22711
rect 14546 22643 14580 22671
rect 14546 22637 14580 22643
rect 14546 22575 14580 22599
rect 14546 22565 14580 22575
rect 14546 22507 14580 22527
rect 14546 22493 14580 22507
rect 14546 22439 14580 22455
rect 14546 22421 14580 22439
rect 14546 22371 14580 22383
rect 14546 22349 14580 22371
rect 14546 22303 14580 22311
rect 14546 22277 14580 22303
rect 14546 22235 14580 22239
rect 14546 22205 14580 22235
rect 14546 22133 14580 22167
rect 14546 22065 14580 22095
rect 14546 22061 14580 22065
rect 14546 21997 14580 22023
rect 14546 21989 14580 21997
rect 14546 21929 14580 21951
rect 14546 21917 14580 21929
rect 14546 21861 14580 21879
rect 14546 21845 14580 21861
rect 14546 21793 14580 21807
rect 14546 21773 14580 21793
rect 14546 21725 14580 21735
rect 14546 21701 14580 21725
rect 14546 21657 14580 21663
rect 14546 21629 14580 21657
rect 14546 21589 14580 21591
rect 14546 21557 14580 21589
rect 14546 21487 14580 21519
rect 14546 21485 14580 21487
rect 14546 21419 14580 21447
rect 14546 21413 14580 21419
rect 14546 21351 14580 21375
rect 14546 21341 14580 21351
rect 14546 21283 14580 21303
rect 14546 21269 14580 21283
rect 14546 21215 14580 21231
rect 14546 21197 14580 21215
rect 14642 23085 14676 23103
rect 14642 23069 14676 23085
rect 14642 23017 14676 23031
rect 14642 22997 14676 23017
rect 14642 22949 14676 22959
rect 14642 22925 14676 22949
rect 14642 22881 14676 22887
rect 14642 22853 14676 22881
rect 14642 22813 14676 22815
rect 14642 22781 14676 22813
rect 14642 22711 14676 22743
rect 14642 22709 14676 22711
rect 14642 22643 14676 22671
rect 14642 22637 14676 22643
rect 14642 22575 14676 22599
rect 14642 22565 14676 22575
rect 14642 22507 14676 22527
rect 14642 22493 14676 22507
rect 14642 22439 14676 22455
rect 14642 22421 14676 22439
rect 14642 22371 14676 22383
rect 14642 22349 14676 22371
rect 14642 22303 14676 22311
rect 14642 22277 14676 22303
rect 14642 22235 14676 22239
rect 14642 22205 14676 22235
rect 14642 22133 14676 22167
rect 14642 22065 14676 22095
rect 14642 22061 14676 22065
rect 14642 21997 14676 22023
rect 14642 21989 14676 21997
rect 14642 21929 14676 21951
rect 14642 21917 14676 21929
rect 14642 21861 14676 21879
rect 14642 21845 14676 21861
rect 14642 21793 14676 21807
rect 14642 21773 14676 21793
rect 14642 21725 14676 21735
rect 14642 21701 14676 21725
rect 14642 21657 14676 21663
rect 14642 21629 14676 21657
rect 14642 21589 14676 21591
rect 14642 21557 14676 21589
rect 14642 21487 14676 21519
rect 14642 21485 14676 21487
rect 14642 21419 14676 21447
rect 14642 21413 14676 21419
rect 14642 21351 14676 21375
rect 14642 21341 14676 21351
rect 14642 21283 14676 21303
rect 14642 21269 14676 21283
rect 14642 21215 14676 21231
rect 14642 21197 14676 21215
rect 14738 23085 14772 23103
rect 14738 23069 14772 23085
rect 14738 23017 14772 23031
rect 14848 23085 14882 23107
rect 14848 23073 14852 23085
rect 14852 23073 14882 23085
rect 14738 22997 14772 23017
rect 14738 22949 14772 22959
rect 14738 22925 14772 22949
rect 14738 22881 14772 22887
rect 14738 22853 14772 22881
rect 14738 22813 14772 22815
rect 14738 22781 14772 22813
rect 14738 22711 14772 22743
rect 14738 22709 14772 22711
rect 14738 22643 14772 22671
rect 14738 22637 14772 22643
rect 14738 22575 14772 22599
rect 14738 22565 14772 22575
rect 14738 22507 14772 22527
rect 14738 22493 14772 22507
rect 14738 22439 14772 22455
rect 14738 22421 14772 22439
rect 14738 22371 14772 22383
rect 14738 22349 14772 22371
rect 14738 22303 14772 22311
rect 14738 22277 14772 22303
rect 14738 22235 14772 22239
rect 14738 22205 14772 22235
rect 14738 22133 14772 22167
rect 14738 22065 14772 22095
rect 14738 22061 14772 22065
rect 14738 21997 14772 22023
rect 14738 21989 14772 21997
rect 14738 21929 14772 21951
rect 14738 21917 14772 21929
rect 14738 21861 14772 21879
rect 14738 21845 14772 21861
rect 14738 21793 14772 21807
rect 14738 21773 14772 21793
rect 14738 21725 14772 21735
rect 14738 21701 14772 21725
rect 14738 21657 14772 21663
rect 14738 21629 14772 21657
rect 14738 21589 14772 21591
rect 14738 21557 14772 21589
rect 14738 21487 14772 21519
rect 14738 21485 14772 21487
rect 14738 21419 14772 21447
rect 14738 21413 14772 21419
rect 14738 21351 14772 21375
rect 14738 21341 14772 21351
rect 14738 21283 14772 21303
rect 14738 21269 14772 21283
rect 14738 21215 14772 21231
rect 14738 21197 14772 21215
rect 14018 21078 14052 21112
rect 14210 21078 14244 21112
rect 14402 21078 14436 21112
rect 14594 21078 14628 21112
rect 15324 23176 15358 23210
rect 15324 23104 15358 23138
rect 15324 23032 15358 23066
rect 15324 22960 15358 22994
rect 15324 22888 15358 22922
rect 15324 22816 15358 22850
rect 15324 21505 15358 21539
rect 15324 21433 15358 21467
rect 15324 21361 15358 21395
rect 15324 21289 15358 21323
rect 15324 21217 15358 21251
rect 15324 21145 15358 21179
rect 15974 23236 16008 23270
rect 15830 23124 15864 23142
rect 15830 23108 15864 23124
rect 15830 23056 15864 23070
rect 15830 23036 15864 23056
rect 15830 22988 15864 22998
rect 15830 22964 15864 22988
rect 15830 22920 15864 22926
rect 15830 22892 15864 22920
rect 15830 22852 15864 22854
rect 15830 22820 15864 22852
rect 15830 22750 15864 22782
rect 15830 22748 15864 22750
rect 15830 22682 15864 22710
rect 15830 22676 15864 22682
rect 15830 22614 15864 22638
rect 15830 22604 15864 22614
rect 15830 22546 15864 22566
rect 15830 22532 15864 22546
rect 15830 22478 15864 22494
rect 15830 22460 15864 22478
rect 15830 22410 15864 22422
rect 15830 22388 15864 22410
rect 15830 22342 15864 22350
rect 15830 22316 15864 22342
rect 15830 22274 15864 22278
rect 15830 22244 15864 22274
rect 15830 22172 15864 22206
rect 15830 22104 15864 22134
rect 15830 22100 15864 22104
rect 15830 22036 15864 22062
rect 15830 22028 15864 22036
rect 15830 21968 15864 21990
rect 15830 21956 15864 21968
rect 15830 21900 15864 21918
rect 15830 21884 15864 21900
rect 15830 21832 15864 21846
rect 15830 21812 15864 21832
rect 15830 21764 15864 21774
rect 15830 21740 15864 21764
rect 15830 21696 15864 21702
rect 15830 21668 15864 21696
rect 15830 21628 15864 21630
rect 15830 21596 15864 21628
rect 15830 21526 15864 21558
rect 15830 21524 15864 21526
rect 15830 21458 15864 21486
rect 15830 21452 15864 21458
rect 15830 21390 15864 21414
rect 15830 21380 15864 21390
rect 15830 21322 15864 21342
rect 15830 21308 15864 21322
rect 15830 21254 15864 21270
rect 15830 21236 15864 21254
rect 15926 23124 15960 23142
rect 15926 23108 15960 23124
rect 15926 23056 15960 23070
rect 15926 23036 15960 23056
rect 15926 22988 15960 22998
rect 15926 22964 15960 22988
rect 15926 22920 15960 22926
rect 15926 22892 15960 22920
rect 15926 22852 15960 22854
rect 15926 22820 15960 22852
rect 15926 22750 15960 22782
rect 15926 22748 15960 22750
rect 15926 22682 15960 22710
rect 15926 22676 15960 22682
rect 15926 22614 15960 22638
rect 15926 22604 15960 22614
rect 15926 22546 15960 22566
rect 15926 22532 15960 22546
rect 15926 22478 15960 22494
rect 15926 22460 15960 22478
rect 15926 22410 15960 22422
rect 15926 22388 15960 22410
rect 15926 22342 15960 22350
rect 15926 22316 15960 22342
rect 15926 22274 15960 22278
rect 15926 22244 15960 22274
rect 15926 22172 15960 22206
rect 15926 22104 15960 22134
rect 15926 22100 15960 22104
rect 15926 22036 15960 22062
rect 15926 22028 15960 22036
rect 15926 21968 15960 21990
rect 15926 21956 15960 21968
rect 15926 21900 15960 21918
rect 15926 21884 15960 21900
rect 15926 21832 15960 21846
rect 15926 21812 15960 21832
rect 15926 21764 15960 21774
rect 15926 21740 15960 21764
rect 15926 21696 15960 21702
rect 15926 21668 15960 21696
rect 15926 21628 15960 21630
rect 15926 21596 15960 21628
rect 15926 21526 15960 21558
rect 15926 21524 15960 21526
rect 15926 21458 15960 21486
rect 15926 21452 15960 21458
rect 15926 21390 15960 21414
rect 15926 21380 15960 21390
rect 15926 21322 15960 21342
rect 15926 21308 15960 21322
rect 15926 21254 15960 21270
rect 15926 21236 15960 21254
rect 16022 23124 16056 23142
rect 16022 23108 16056 23124
rect 16022 23056 16056 23070
rect 16022 23036 16056 23056
rect 16022 22988 16056 22998
rect 16022 22964 16056 22988
rect 16022 22920 16056 22926
rect 16022 22892 16056 22920
rect 16022 22852 16056 22854
rect 16022 22820 16056 22852
rect 16022 22750 16056 22782
rect 16022 22748 16056 22750
rect 16022 22682 16056 22710
rect 16022 22676 16056 22682
rect 16022 22614 16056 22638
rect 16022 22604 16056 22614
rect 16022 22546 16056 22566
rect 16022 22532 16056 22546
rect 16022 22478 16056 22494
rect 16022 22460 16056 22478
rect 16022 22410 16056 22422
rect 16022 22388 16056 22410
rect 16022 22342 16056 22350
rect 16022 22316 16056 22342
rect 16022 22274 16056 22278
rect 16022 22244 16056 22274
rect 16022 22172 16056 22206
rect 16022 22104 16056 22134
rect 16022 22100 16056 22104
rect 16022 22036 16056 22062
rect 16022 22028 16056 22036
rect 16022 21968 16056 21990
rect 16022 21956 16056 21968
rect 16022 21900 16056 21918
rect 16022 21884 16056 21900
rect 16022 21832 16056 21846
rect 16022 21812 16056 21832
rect 16022 21764 16056 21774
rect 16022 21740 16056 21764
rect 16022 21696 16056 21702
rect 16022 21668 16056 21696
rect 16022 21628 16056 21630
rect 16022 21596 16056 21628
rect 16022 21526 16056 21558
rect 16022 21524 16056 21526
rect 16022 21458 16056 21486
rect 16022 21452 16056 21458
rect 16022 21390 16056 21414
rect 16022 21380 16056 21390
rect 16022 21322 16056 21342
rect 16022 21308 16056 21322
rect 16022 21254 16056 21270
rect 16022 21236 16056 21254
rect 16118 23124 16152 23142
rect 16118 23108 16152 23124
rect 16118 23056 16152 23070
rect 16118 23036 16152 23056
rect 16118 22988 16152 22998
rect 16118 22964 16152 22988
rect 16118 22920 16152 22926
rect 16118 22892 16152 22920
rect 16118 22852 16152 22854
rect 16118 22820 16152 22852
rect 16118 22750 16152 22782
rect 16118 22748 16152 22750
rect 16118 22682 16152 22710
rect 16118 22676 16152 22682
rect 16118 22614 16152 22638
rect 16118 22604 16152 22614
rect 16118 22546 16152 22566
rect 16118 22532 16152 22546
rect 16118 22478 16152 22494
rect 16118 22460 16152 22478
rect 16118 22410 16152 22422
rect 16118 22388 16152 22410
rect 16118 22342 16152 22350
rect 16118 22316 16152 22342
rect 16118 22274 16152 22278
rect 16118 22244 16152 22274
rect 16118 22172 16152 22206
rect 16118 22104 16152 22134
rect 16118 22100 16152 22104
rect 16118 22036 16152 22062
rect 16118 22028 16152 22036
rect 16118 21968 16152 21990
rect 16118 21956 16152 21968
rect 16118 21900 16152 21918
rect 16118 21884 16152 21900
rect 16118 21832 16152 21846
rect 16118 21812 16152 21832
rect 16662 23975 16696 23993
rect 16662 23959 16696 23975
rect 16662 23907 16696 23921
rect 16662 23887 16696 23907
rect 16662 23839 16696 23849
rect 16662 23815 16696 23839
rect 16662 23771 16696 23777
rect 16662 23743 16696 23771
rect 16662 23703 16696 23705
rect 16662 23671 16696 23703
rect 16662 23601 16696 23633
rect 16662 23599 16696 23601
rect 16662 23533 16696 23561
rect 16662 23527 16696 23533
rect 16662 23465 16696 23489
rect 16662 23455 16696 23465
rect 16662 23397 16696 23417
rect 16662 23383 16696 23397
rect 16662 23329 16696 23345
rect 16662 23311 16696 23329
rect 16662 23261 16696 23273
rect 16662 23239 16696 23261
rect 16662 23193 16696 23201
rect 16662 23167 16696 23193
rect 16662 23125 16696 23129
rect 16662 23095 16696 23125
rect 16662 23023 16696 23057
rect 16662 22955 16696 22985
rect 16662 22951 16696 22955
rect 16662 22887 16696 22913
rect 16662 22879 16696 22887
rect 16662 22819 16696 22841
rect 16662 22807 16696 22819
rect 16662 22751 16696 22769
rect 16662 22735 16696 22751
rect 16662 22683 16696 22697
rect 16662 22663 16696 22683
rect 16662 22615 16696 22625
rect 16662 22591 16696 22615
rect 16662 22547 16696 22553
rect 16662 22519 16696 22547
rect 16662 22479 16696 22481
rect 16662 22447 16696 22479
rect 16662 22377 16696 22409
rect 16662 22375 16696 22377
rect 16662 22309 16696 22337
rect 16662 22303 16696 22309
rect 16662 22241 16696 22265
rect 16662 22231 16696 22241
rect 16662 22173 16696 22193
rect 16662 22159 16696 22173
rect 16662 22105 16696 22121
rect 16662 22087 16696 22105
rect 16758 23975 16792 23993
rect 16758 23959 16792 23975
rect 16758 23907 16792 23921
rect 16758 23887 16792 23907
rect 16758 23839 16792 23849
rect 16758 23815 16792 23839
rect 16758 23771 16792 23777
rect 16758 23743 16792 23771
rect 16758 23703 16792 23705
rect 16758 23671 16792 23703
rect 16758 23601 16792 23633
rect 16758 23599 16792 23601
rect 16758 23533 16792 23561
rect 16758 23527 16792 23533
rect 16758 23465 16792 23489
rect 16758 23455 16792 23465
rect 16758 23397 16792 23417
rect 16758 23383 16792 23397
rect 16758 23329 16792 23345
rect 16758 23311 16792 23329
rect 16758 23261 16792 23273
rect 16758 23239 16792 23261
rect 16758 23193 16792 23201
rect 16758 23167 16792 23193
rect 16758 23125 16792 23129
rect 16758 23095 16792 23125
rect 16758 23023 16792 23057
rect 16758 22955 16792 22985
rect 16758 22951 16792 22955
rect 16758 22887 16792 22913
rect 16758 22879 16792 22887
rect 16758 22819 16792 22841
rect 16758 22807 16792 22819
rect 16758 22751 16792 22769
rect 16758 22735 16792 22751
rect 16758 22683 16792 22697
rect 16758 22663 16792 22683
rect 16758 22615 16792 22625
rect 16758 22591 16792 22615
rect 16758 22547 16792 22553
rect 16758 22519 16792 22547
rect 16758 22479 16792 22481
rect 16758 22447 16792 22479
rect 16758 22377 16792 22409
rect 16758 22375 16792 22377
rect 16758 22309 16792 22337
rect 16758 22303 16792 22309
rect 16758 22241 16792 22265
rect 16758 22231 16792 22241
rect 16758 22173 16792 22193
rect 16758 22159 16792 22173
rect 16758 22105 16792 22121
rect 16758 22087 16792 22105
rect 16854 23975 16888 23993
rect 16854 23959 16888 23975
rect 16854 23907 16888 23921
rect 16854 23887 16888 23907
rect 16854 23839 16888 23849
rect 16854 23815 16888 23839
rect 16854 23771 16888 23777
rect 16854 23743 16888 23771
rect 16854 23703 16888 23705
rect 16854 23671 16888 23703
rect 16854 23601 16888 23633
rect 16854 23599 16888 23601
rect 16854 23533 16888 23561
rect 16854 23527 16888 23533
rect 16854 23465 16888 23489
rect 16854 23455 16888 23465
rect 16854 23397 16888 23417
rect 16854 23383 16888 23397
rect 16854 23329 16888 23345
rect 16854 23311 16888 23329
rect 16854 23261 16888 23273
rect 16854 23239 16888 23261
rect 16854 23193 16888 23201
rect 16854 23167 16888 23193
rect 16854 23125 16888 23129
rect 16854 23095 16888 23125
rect 16854 23023 16888 23057
rect 16854 22955 16888 22985
rect 16854 22951 16888 22955
rect 16854 22887 16888 22913
rect 16854 22879 16888 22887
rect 16854 22819 16888 22841
rect 16854 22807 16888 22819
rect 16854 22751 16888 22769
rect 16854 22735 16888 22751
rect 16854 22683 16888 22697
rect 16854 22663 16888 22683
rect 16854 22615 16888 22625
rect 16854 22591 16888 22615
rect 16854 22547 16888 22553
rect 16854 22519 16888 22547
rect 16854 22479 16888 22481
rect 16854 22447 16888 22479
rect 16854 22377 16888 22409
rect 16854 22375 16888 22377
rect 16854 22309 16888 22337
rect 16854 22303 16888 22309
rect 16854 22241 16888 22265
rect 16854 22231 16888 22241
rect 16854 22173 16888 22193
rect 16854 22159 16888 22173
rect 16854 22105 16888 22121
rect 16854 22087 16888 22105
rect 16950 23975 16984 23993
rect 16950 23959 16984 23975
rect 16950 23907 16984 23921
rect 16950 23887 16984 23907
rect 16950 23839 16984 23849
rect 16950 23815 16984 23839
rect 16950 23771 16984 23777
rect 16950 23743 16984 23771
rect 16950 23703 16984 23705
rect 16950 23671 16984 23703
rect 16950 23601 16984 23633
rect 16950 23599 16984 23601
rect 16950 23533 16984 23561
rect 16950 23527 16984 23533
rect 16950 23465 16984 23489
rect 16950 23455 16984 23465
rect 16950 23397 16984 23417
rect 16950 23383 16984 23397
rect 16950 23329 16984 23345
rect 16950 23311 16984 23329
rect 16950 23261 16984 23273
rect 16950 23239 16984 23261
rect 16950 23193 16984 23201
rect 16950 23167 16984 23193
rect 16950 23125 16984 23129
rect 16950 23095 16984 23125
rect 16950 23023 16984 23057
rect 16950 22955 16984 22985
rect 16950 22951 16984 22955
rect 16950 22887 16984 22913
rect 16950 22879 16984 22887
rect 16950 22819 16984 22841
rect 16950 22807 16984 22819
rect 16950 22751 16984 22769
rect 16950 22735 16984 22751
rect 16950 22683 16984 22697
rect 16950 22663 16984 22683
rect 16950 22615 16984 22625
rect 16950 22591 16984 22615
rect 16950 22547 16984 22553
rect 16950 22519 16984 22547
rect 16950 22479 16984 22481
rect 16950 22447 16984 22479
rect 16950 22377 16984 22409
rect 16950 22375 16984 22377
rect 16950 22309 16984 22337
rect 16950 22303 16984 22309
rect 16950 22241 16984 22265
rect 16950 22231 16984 22241
rect 16950 22173 16984 22193
rect 16950 22159 16984 22173
rect 16950 22105 16984 22121
rect 16950 22087 16984 22105
rect 17046 23975 17080 23993
rect 17046 23959 17080 23975
rect 17046 23907 17080 23921
rect 17046 23887 17080 23907
rect 17046 23839 17080 23849
rect 17046 23815 17080 23839
rect 17046 23771 17080 23777
rect 17046 23743 17080 23771
rect 17046 23703 17080 23705
rect 17046 23671 17080 23703
rect 17046 23601 17080 23633
rect 17046 23599 17080 23601
rect 17046 23533 17080 23561
rect 17046 23527 17080 23533
rect 17046 23465 17080 23489
rect 17046 23455 17080 23465
rect 17046 23397 17080 23417
rect 17046 23383 17080 23397
rect 17046 23329 17080 23345
rect 17046 23311 17080 23329
rect 17046 23261 17080 23273
rect 17046 23239 17080 23261
rect 17046 23193 17080 23201
rect 17046 23167 17080 23193
rect 17046 23125 17080 23129
rect 17046 23095 17080 23125
rect 17046 23023 17080 23057
rect 17046 22955 17080 22985
rect 17046 22951 17080 22955
rect 17046 22887 17080 22913
rect 17046 22879 17080 22887
rect 17046 22819 17080 22841
rect 17046 22807 17080 22819
rect 17046 22751 17080 22769
rect 17046 22735 17080 22751
rect 17046 22683 17080 22697
rect 17046 22663 17080 22683
rect 17046 22615 17080 22625
rect 17046 22591 17080 22615
rect 17046 22547 17080 22553
rect 17046 22519 17080 22547
rect 17046 22479 17080 22481
rect 17046 22447 17080 22479
rect 17046 22377 17080 22409
rect 17046 22375 17080 22377
rect 17046 22309 17080 22337
rect 17046 22303 17080 22309
rect 17046 22241 17080 22265
rect 17046 22231 17080 22241
rect 17046 22173 17080 22193
rect 17046 22159 17080 22173
rect 17046 22105 17080 22121
rect 17046 22087 17080 22105
rect 17142 23975 17176 23993
rect 17142 23959 17176 23975
rect 17142 23907 17176 23921
rect 17142 23887 17176 23907
rect 17142 23839 17176 23849
rect 17142 23815 17176 23839
rect 17142 23771 17176 23777
rect 17142 23743 17176 23771
rect 17142 23703 17176 23705
rect 17142 23671 17176 23703
rect 17142 23601 17176 23633
rect 17142 23599 17176 23601
rect 17142 23533 17176 23561
rect 17142 23527 17176 23533
rect 17142 23465 17176 23489
rect 17142 23455 17176 23465
rect 17142 23397 17176 23417
rect 17142 23383 17176 23397
rect 17142 23329 17176 23345
rect 17142 23311 17176 23329
rect 17142 23261 17176 23273
rect 17142 23239 17176 23261
rect 17142 23193 17176 23201
rect 17142 23167 17176 23193
rect 17142 23125 17176 23129
rect 17142 23095 17176 23125
rect 17142 23023 17176 23057
rect 17142 22955 17176 22985
rect 17142 22951 17176 22955
rect 17142 22887 17176 22913
rect 17142 22879 17176 22887
rect 17142 22819 17176 22841
rect 17142 22807 17176 22819
rect 17142 22751 17176 22769
rect 17142 22735 17176 22751
rect 17142 22683 17176 22697
rect 17142 22663 17176 22683
rect 17142 22615 17176 22625
rect 17142 22591 17176 22615
rect 17142 22547 17176 22553
rect 17142 22519 17176 22547
rect 17142 22479 17176 22481
rect 17142 22447 17176 22479
rect 17142 22377 17176 22409
rect 17142 22375 17176 22377
rect 17142 22309 17176 22337
rect 17142 22303 17176 22309
rect 17142 22241 17176 22265
rect 17142 22231 17176 22241
rect 17142 22173 17176 22193
rect 17142 22159 17176 22173
rect 17142 22105 17176 22121
rect 17142 22087 17176 22105
rect 17238 23975 17272 23993
rect 17238 23959 17272 23975
rect 17238 23907 17272 23921
rect 17238 23887 17272 23907
rect 17238 23839 17272 23849
rect 17238 23815 17272 23839
rect 17238 23771 17272 23777
rect 17238 23743 17272 23771
rect 17238 23703 17272 23705
rect 17238 23671 17272 23703
rect 17238 23601 17272 23633
rect 17238 23599 17272 23601
rect 17238 23533 17272 23561
rect 17238 23527 17272 23533
rect 17238 23465 17272 23489
rect 17238 23455 17272 23465
rect 17238 23397 17272 23417
rect 17238 23383 17272 23397
rect 17238 23329 17272 23345
rect 17238 23311 17272 23329
rect 17238 23261 17272 23273
rect 17238 23239 17272 23261
rect 17238 23193 17272 23201
rect 17238 23167 17272 23193
rect 17238 23125 17272 23129
rect 17238 23095 17272 23125
rect 17238 23023 17272 23057
rect 17238 22955 17272 22985
rect 17238 22951 17272 22955
rect 17238 22887 17272 22913
rect 17238 22879 17272 22887
rect 17238 22819 17272 22841
rect 17238 22807 17272 22819
rect 17238 22751 17272 22769
rect 17238 22735 17272 22751
rect 17238 22683 17272 22697
rect 17238 22663 17272 22683
rect 17238 22615 17272 22625
rect 17238 22591 17272 22615
rect 17238 22547 17272 22553
rect 17238 22519 17272 22547
rect 17238 22479 17272 22481
rect 17238 22447 17272 22479
rect 17238 22377 17272 22409
rect 17238 22375 17272 22377
rect 17238 22309 17272 22337
rect 17238 22303 17272 22309
rect 17238 22241 17272 22265
rect 17238 22231 17272 22241
rect 17238 22173 17272 22193
rect 17238 22159 17272 22173
rect 17238 22105 17272 22121
rect 17238 22087 17272 22105
rect 17334 23975 17368 23993
rect 17334 23959 17368 23975
rect 17334 23907 17368 23921
rect 17334 23887 17368 23907
rect 17334 23839 17368 23849
rect 17334 23815 17368 23839
rect 17334 23771 17368 23777
rect 17334 23743 17368 23771
rect 17334 23703 17368 23705
rect 17334 23671 17368 23703
rect 17334 23601 17368 23633
rect 17334 23599 17368 23601
rect 17334 23533 17368 23561
rect 17334 23527 17368 23533
rect 17334 23465 17368 23489
rect 17334 23455 17368 23465
rect 17334 23397 17368 23417
rect 17334 23383 17368 23397
rect 17334 23329 17368 23345
rect 17334 23311 17368 23329
rect 17334 23261 17368 23273
rect 17334 23239 17368 23261
rect 17334 23193 17368 23201
rect 17334 23167 17368 23193
rect 17334 23125 17368 23129
rect 17334 23095 17368 23125
rect 17334 23023 17368 23057
rect 17334 22955 17368 22985
rect 17334 22951 17368 22955
rect 17334 22887 17368 22913
rect 17334 22879 17368 22887
rect 17334 22819 17368 22841
rect 17334 22807 17368 22819
rect 17334 22751 17368 22769
rect 17334 22735 17368 22751
rect 17334 22683 17368 22697
rect 17334 22663 17368 22683
rect 17334 22615 17368 22625
rect 17334 22591 17368 22615
rect 17334 22547 17368 22553
rect 17334 22519 17368 22547
rect 17334 22479 17368 22481
rect 17334 22447 17368 22479
rect 17334 22377 17368 22409
rect 17334 22375 17368 22377
rect 17334 22309 17368 22337
rect 17334 22303 17368 22309
rect 17334 22241 17368 22265
rect 17334 22231 17368 22241
rect 17334 22173 17368 22193
rect 17334 22159 17368 22173
rect 17334 22105 17368 22121
rect 17334 22087 17368 22105
rect 17430 23975 17464 23993
rect 17430 23959 17464 23975
rect 17430 23907 17464 23921
rect 17430 23887 17464 23907
rect 17430 23839 17464 23849
rect 17430 23815 17464 23839
rect 17430 23771 17464 23777
rect 17430 23743 17464 23771
rect 17430 23703 17464 23705
rect 17430 23671 17464 23703
rect 17430 23601 17464 23633
rect 17430 23599 17464 23601
rect 17430 23533 17464 23561
rect 17430 23527 17464 23533
rect 17430 23465 17464 23489
rect 17430 23455 17464 23465
rect 17430 23397 17464 23417
rect 17430 23383 17464 23397
rect 17430 23329 17464 23345
rect 17430 23311 17464 23329
rect 17430 23261 17464 23273
rect 17430 23239 17464 23261
rect 17430 23193 17464 23201
rect 17430 23167 17464 23193
rect 17430 23125 17464 23129
rect 17430 23095 17464 23125
rect 17430 23023 17464 23057
rect 17430 22955 17464 22985
rect 17430 22951 17464 22955
rect 17430 22887 17464 22913
rect 17430 22879 17464 22887
rect 17430 22819 17464 22841
rect 17430 22807 17464 22819
rect 17430 22751 17464 22769
rect 17430 22735 17464 22751
rect 17430 22683 17464 22697
rect 17430 22663 17464 22683
rect 17430 22615 17464 22625
rect 17430 22591 17464 22615
rect 17430 22547 17464 22553
rect 17430 22519 17464 22547
rect 17430 22479 17464 22481
rect 17430 22447 17464 22479
rect 17430 22377 17464 22409
rect 17430 22375 17464 22377
rect 17430 22309 17464 22337
rect 17430 22303 17464 22309
rect 17430 22241 17464 22265
rect 17430 22231 17464 22241
rect 17430 22173 17464 22193
rect 17430 22159 17464 22173
rect 17430 22105 17464 22121
rect 17430 22087 17464 22105
rect 17526 23975 17560 23993
rect 17526 23959 17560 23975
rect 17526 23907 17560 23921
rect 17526 23887 17560 23907
rect 17526 23839 17560 23849
rect 17526 23815 17560 23839
rect 17526 23771 17560 23777
rect 17526 23743 17560 23771
rect 17526 23703 17560 23705
rect 17526 23671 17560 23703
rect 17526 23601 17560 23633
rect 17526 23599 17560 23601
rect 17526 23533 17560 23561
rect 17526 23527 17560 23533
rect 17526 23465 17560 23489
rect 17526 23455 17560 23465
rect 17526 23397 17560 23417
rect 17526 23383 17560 23397
rect 17526 23329 17560 23345
rect 17526 23311 17560 23329
rect 17526 23261 17560 23273
rect 17526 23239 17560 23261
rect 17526 23193 17560 23201
rect 17526 23167 17560 23193
rect 17526 23125 17560 23129
rect 17526 23095 17560 23125
rect 17526 23023 17560 23057
rect 17526 22955 17560 22985
rect 17526 22951 17560 22955
rect 17526 22887 17560 22913
rect 17526 22879 17560 22887
rect 17526 22819 17560 22841
rect 17526 22807 17560 22819
rect 17526 22751 17560 22769
rect 17526 22735 17560 22751
rect 17526 22683 17560 22697
rect 17526 22663 17560 22683
rect 17526 22615 17560 22625
rect 17526 22591 17560 22615
rect 17526 22547 17560 22553
rect 17526 22519 17560 22547
rect 17526 22479 17560 22481
rect 17526 22447 17560 22479
rect 17526 22377 17560 22409
rect 17526 22375 17560 22377
rect 17526 22309 17560 22337
rect 17526 22303 17560 22309
rect 17526 22241 17560 22265
rect 17526 22231 17560 22241
rect 17526 22173 17560 22193
rect 17526 22159 17560 22173
rect 17526 22105 17560 22121
rect 17526 22087 17560 22105
rect 17622 23975 17656 23993
rect 17622 23959 17656 23975
rect 17622 23907 17656 23921
rect 17622 23887 17656 23907
rect 17622 23839 17656 23849
rect 17622 23815 17656 23839
rect 17622 23771 17656 23777
rect 17622 23743 17656 23771
rect 17622 23703 17656 23705
rect 17622 23671 17656 23703
rect 17622 23601 17656 23633
rect 17622 23599 17656 23601
rect 17622 23533 17656 23561
rect 17622 23527 17656 23533
rect 17622 23465 17656 23489
rect 17622 23455 17656 23465
rect 17622 23397 17656 23417
rect 17622 23383 17656 23397
rect 17622 23329 17656 23345
rect 17622 23311 17656 23329
rect 17622 23261 17656 23273
rect 17622 23239 17656 23261
rect 17622 23193 17656 23201
rect 17622 23167 17656 23193
rect 17622 23125 17656 23129
rect 17622 23095 17656 23125
rect 17622 23023 17656 23057
rect 17622 22955 17656 22985
rect 17622 22951 17656 22955
rect 17622 22887 17656 22913
rect 17622 22879 17656 22887
rect 17622 22819 17656 22841
rect 17622 22807 17656 22819
rect 17622 22751 17656 22769
rect 17622 22735 17656 22751
rect 17622 22683 17656 22697
rect 17622 22663 17656 22683
rect 17622 22615 17656 22625
rect 17622 22591 17656 22615
rect 17622 22547 17656 22553
rect 17622 22519 17656 22547
rect 17622 22479 17656 22481
rect 17622 22447 17656 22479
rect 17622 22377 17656 22409
rect 17622 22375 17656 22377
rect 17622 22309 17656 22337
rect 17622 22303 17656 22309
rect 17622 22241 17656 22265
rect 17622 22231 17656 22241
rect 17622 22173 17656 22193
rect 17622 22159 17656 22173
rect 17622 22105 17656 22121
rect 17622 22087 17656 22105
rect 16710 21968 16744 22002
rect 16902 21968 16936 22002
rect 17094 21968 17128 22002
rect 17286 21968 17320 22002
rect 17478 21968 17512 22002
rect 16118 21764 16152 21774
rect 16118 21740 16152 21764
rect 16118 21696 16152 21702
rect 16118 21668 16152 21696
rect 16118 21628 16152 21630
rect 16118 21596 16152 21628
rect 17387 21612 17493 21718
rect 16118 21526 16152 21558
rect 16118 21524 16152 21526
rect 16118 21458 16152 21486
rect 16118 21452 16152 21458
rect 16118 21390 16152 21414
rect 16118 21380 16152 21390
rect 16118 21322 16152 21342
rect 16118 21308 16152 21322
rect 16118 21254 16152 21270
rect 16118 21236 16152 21254
rect 15878 21108 15912 21142
rect 16070 21108 16104 21142
rect 16804 21296 16838 21330
rect 16804 21224 16838 21258
rect 16804 21152 16838 21186
rect 16804 21080 16838 21114
rect 16804 21008 16838 21042
rect 16804 20936 16838 20970
rect 14974 20484 15008 20518
rect 15166 20484 15200 20518
rect 15358 20484 15392 20518
rect 13331 19608 13725 19714
rect 13900 19608 14294 19714
rect 13331 19222 13725 19328
rect 13900 19222 14294 19328
rect 14830 20398 14864 20432
rect 14830 20330 14864 20360
rect 14830 20326 14864 20330
rect 14830 20262 14864 20288
rect 14830 20254 14864 20262
rect 14830 20194 14864 20216
rect 14830 20182 14864 20194
rect 14830 20126 14864 20144
rect 14830 20110 14864 20126
rect 14830 20058 14864 20072
rect 14830 20038 14864 20058
rect 14830 19990 14864 20000
rect 14830 19966 14864 19990
rect 14830 19922 14864 19928
rect 14830 19894 14864 19922
rect 14830 19854 14864 19856
rect 14830 19822 14864 19854
rect 14830 19752 14864 19784
rect 14830 19750 14864 19752
rect 14830 19684 14864 19712
rect 14830 19678 14864 19684
rect 14830 19616 14864 19640
rect 14830 19606 14864 19616
rect 14830 19548 14864 19568
rect 14830 19534 14864 19548
rect 14830 19480 14864 19496
rect 14830 19462 14864 19480
rect 14830 19412 14864 19424
rect 14830 19390 14864 19412
rect 14830 19344 14864 19352
rect 14830 19318 14864 19344
rect 14926 20398 14960 20432
rect 14926 20330 14960 20360
rect 14926 20326 14960 20330
rect 14926 20262 14960 20288
rect 14926 20254 14960 20262
rect 14926 20194 14960 20216
rect 14926 20182 14960 20194
rect 14926 20126 14960 20144
rect 14926 20110 14960 20126
rect 14926 20058 14960 20072
rect 14926 20038 14960 20058
rect 14926 19990 14960 20000
rect 14926 19966 14960 19990
rect 14926 19922 14960 19928
rect 14926 19894 14960 19922
rect 14926 19854 14960 19856
rect 14926 19822 14960 19854
rect 14926 19752 14960 19784
rect 14926 19750 14960 19752
rect 14926 19684 14960 19712
rect 14926 19678 14960 19684
rect 14926 19616 14960 19640
rect 14926 19606 14960 19616
rect 14926 19548 14960 19568
rect 14926 19534 14960 19548
rect 14926 19480 14960 19496
rect 14926 19462 14960 19480
rect 14926 19412 14960 19424
rect 14926 19390 14960 19412
rect 14926 19344 14960 19352
rect 14926 19318 14960 19344
rect 14830 19276 14864 19280
rect 14830 19246 14864 19276
rect 14830 19174 14864 19208
rect 14926 19276 14960 19280
rect 14926 19246 14960 19276
rect 14926 19174 14960 19208
rect 15022 20398 15056 20432
rect 15022 20330 15056 20360
rect 15022 20326 15056 20330
rect 15022 20262 15056 20288
rect 15022 20254 15056 20262
rect 15022 20194 15056 20216
rect 15022 20182 15056 20194
rect 15022 20126 15056 20144
rect 15022 20110 15056 20126
rect 15022 20058 15056 20072
rect 15022 20038 15056 20058
rect 15022 19990 15056 20000
rect 15022 19966 15056 19990
rect 15022 19922 15056 19928
rect 15022 19894 15056 19922
rect 15022 19854 15056 19856
rect 15022 19822 15056 19854
rect 15022 19752 15056 19784
rect 15022 19750 15056 19752
rect 15022 19684 15056 19712
rect 15022 19678 15056 19684
rect 15022 19616 15056 19640
rect 15022 19606 15056 19616
rect 15022 19548 15056 19568
rect 15022 19534 15056 19548
rect 15022 19480 15056 19496
rect 15022 19462 15056 19480
rect 15022 19412 15056 19424
rect 15022 19390 15056 19412
rect 15022 19344 15056 19352
rect 15022 19318 15056 19344
rect 15022 19276 15056 19280
rect 15022 19246 15056 19276
rect 15022 19174 15056 19208
rect 15118 20398 15152 20432
rect 15118 20330 15152 20360
rect 15118 20326 15152 20330
rect 15118 20262 15152 20288
rect 15118 20254 15152 20262
rect 15118 20194 15152 20216
rect 15118 20182 15152 20194
rect 15118 20126 15152 20144
rect 15118 20110 15152 20126
rect 15118 20058 15152 20072
rect 15118 20038 15152 20058
rect 15118 19990 15152 20000
rect 15118 19966 15152 19990
rect 15118 19922 15152 19928
rect 15118 19894 15152 19922
rect 15118 19854 15152 19856
rect 15118 19822 15152 19854
rect 15118 19752 15152 19784
rect 15118 19750 15152 19752
rect 15118 19684 15152 19712
rect 15118 19678 15152 19684
rect 15118 19616 15152 19640
rect 15118 19606 15152 19616
rect 15118 19548 15152 19568
rect 15118 19534 15152 19548
rect 15118 19480 15152 19496
rect 15118 19462 15152 19480
rect 15118 19412 15152 19424
rect 15118 19390 15152 19412
rect 15118 19344 15152 19352
rect 15118 19318 15152 19344
rect 15118 19276 15152 19280
rect 15118 19246 15152 19276
rect 15118 19174 15152 19208
rect 15214 20398 15248 20432
rect 15214 20330 15248 20360
rect 15214 20326 15248 20330
rect 15214 20262 15248 20288
rect 15214 20254 15248 20262
rect 15214 20194 15248 20216
rect 15214 20182 15248 20194
rect 15214 20126 15248 20144
rect 15214 20110 15248 20126
rect 15214 20058 15248 20072
rect 15214 20038 15248 20058
rect 15214 19990 15248 20000
rect 15214 19966 15248 19990
rect 15214 19922 15248 19928
rect 15214 19894 15248 19922
rect 15214 19854 15248 19856
rect 15214 19822 15248 19854
rect 15214 19752 15248 19784
rect 15214 19750 15248 19752
rect 15214 19684 15248 19712
rect 15214 19678 15248 19684
rect 15214 19616 15248 19640
rect 15214 19606 15248 19616
rect 15214 19548 15248 19568
rect 15214 19534 15248 19548
rect 15214 19480 15248 19496
rect 15214 19462 15248 19480
rect 15214 19412 15248 19424
rect 15214 19390 15248 19412
rect 15214 19344 15248 19352
rect 15214 19318 15248 19344
rect 15214 19276 15248 19280
rect 15214 19246 15248 19276
rect 15214 19174 15248 19208
rect 15310 20398 15344 20432
rect 15310 20330 15344 20360
rect 15310 20326 15344 20330
rect 15310 20262 15344 20288
rect 15310 20254 15344 20262
rect 15310 20194 15344 20216
rect 15310 20182 15344 20194
rect 15310 20126 15344 20144
rect 15310 20110 15344 20126
rect 15310 20058 15344 20072
rect 15310 20038 15344 20058
rect 15310 19990 15344 20000
rect 15310 19966 15344 19990
rect 15310 19922 15344 19928
rect 15310 19894 15344 19922
rect 15310 19854 15344 19856
rect 15310 19822 15344 19854
rect 15310 19752 15344 19784
rect 15310 19750 15344 19752
rect 15310 19684 15344 19712
rect 15310 19678 15344 19684
rect 15310 19616 15344 19640
rect 15310 19606 15344 19616
rect 15310 19548 15344 19568
rect 15310 19534 15344 19548
rect 15310 19480 15344 19496
rect 15310 19462 15344 19480
rect 15310 19412 15344 19424
rect 15310 19390 15344 19412
rect 15310 19344 15344 19352
rect 15310 19318 15344 19344
rect 15310 19276 15344 19280
rect 15310 19246 15344 19276
rect 15310 19174 15344 19208
rect 15406 20398 15440 20432
rect 15406 20330 15440 20360
rect 15406 20326 15440 20330
rect 15406 20262 15440 20288
rect 15406 20254 15440 20262
rect 15406 20194 15440 20216
rect 15406 20182 15440 20194
rect 15406 20126 15440 20144
rect 15406 20110 15440 20126
rect 15406 20058 15440 20072
rect 15406 20038 15440 20058
rect 15406 19990 15440 20000
rect 15406 19966 15440 19990
rect 15406 19922 15440 19928
rect 15406 19894 15440 19922
rect 15406 19854 15440 19856
rect 15406 19822 15440 19854
rect 15406 19752 15440 19784
rect 15406 19750 15440 19752
rect 15406 19684 15440 19712
rect 15406 19678 15440 19684
rect 15406 19616 15440 19640
rect 15406 19606 15440 19616
rect 15406 19548 15440 19568
rect 15406 19534 15440 19548
rect 15406 19480 15440 19496
rect 15406 19462 15440 19480
rect 15406 19412 15440 19424
rect 15406 19390 15440 19412
rect 15406 19344 15440 19352
rect 15406 19318 15440 19344
rect 15406 19276 15440 19280
rect 15406 19246 15440 19276
rect 15406 19174 15440 19208
rect 15502 20398 15536 20432
rect 15502 20330 15536 20360
rect 15502 20326 15536 20330
rect 15502 20262 15536 20288
rect 15502 20254 15536 20262
rect 15502 20194 15536 20216
rect 15502 20182 15536 20194
rect 15502 20126 15536 20144
rect 15502 20110 15536 20126
rect 15502 20058 15536 20072
rect 15502 20038 15536 20058
rect 15502 19990 15536 20000
rect 15502 19966 15536 19990
rect 15502 19922 15536 19928
rect 15502 19894 15536 19922
rect 15502 19854 15536 19856
rect 15502 19822 15536 19854
rect 15502 19752 15536 19784
rect 15502 19750 15536 19752
rect 15502 19684 15536 19712
rect 15502 19678 15536 19684
rect 15502 19616 15536 19640
rect 15502 19606 15536 19616
rect 15502 19548 15536 19568
rect 15502 19534 15536 19548
rect 15502 19480 15536 19496
rect 15502 19462 15536 19480
rect 15502 19412 15536 19424
rect 15502 19390 15536 19412
rect 15502 19344 15536 19352
rect 15502 19318 15536 19344
rect 15502 19276 15536 19280
rect 15502 19246 15536 19276
rect 15502 19174 15536 19208
rect 14878 19088 14912 19122
rect 15070 19088 15104 19122
rect 15262 19088 15296 19122
rect 15454 19088 15488 19122
rect 16134 19998 16168 20032
rect 15990 19917 16024 19937
rect 15990 19903 16024 19917
rect 15990 19849 16024 19865
rect 15990 19831 16024 19849
rect 15990 19781 16024 19793
rect 15990 19759 16024 19781
rect 15990 19713 16024 19721
rect 15990 19687 16024 19713
rect 15990 19645 16024 19649
rect 15990 19615 16024 19645
rect 15990 19543 16024 19577
rect 15990 19475 16024 19505
rect 15990 19471 16024 19475
rect 15990 19407 16024 19433
rect 15990 19399 16024 19407
rect 15990 19339 16024 19361
rect 15990 19327 16024 19339
rect 15990 19271 16024 19289
rect 15990 19255 16024 19271
rect 15990 19203 16024 19217
rect 15990 19183 16024 19203
rect 16086 19917 16120 19937
rect 16086 19903 16120 19917
rect 16086 19849 16120 19865
rect 16086 19831 16120 19849
rect 16086 19781 16120 19793
rect 16086 19759 16120 19781
rect 16086 19713 16120 19721
rect 16086 19687 16120 19713
rect 16086 19645 16120 19649
rect 16086 19615 16120 19645
rect 16086 19543 16120 19577
rect 16086 19475 16120 19505
rect 16086 19471 16120 19475
rect 16086 19407 16120 19433
rect 16086 19399 16120 19407
rect 16086 19339 16120 19361
rect 16086 19327 16120 19339
rect 16086 19271 16120 19289
rect 16086 19255 16120 19271
rect 16086 19203 16120 19217
rect 16086 19183 16120 19203
rect 16182 19917 16216 19937
rect 16182 19903 16216 19917
rect 16182 19849 16216 19865
rect 16182 19831 16216 19849
rect 16182 19781 16216 19793
rect 16182 19759 16216 19781
rect 16182 19713 16216 19721
rect 16182 19687 16216 19713
rect 16182 19645 16216 19649
rect 16182 19615 16216 19645
rect 16182 19543 16216 19577
rect 16182 19475 16216 19505
rect 16182 19471 16216 19475
rect 16182 19407 16216 19433
rect 16182 19399 16216 19407
rect 16182 19339 16216 19361
rect 16182 19327 16216 19339
rect 16182 19271 16216 19289
rect 16182 19255 16216 19271
rect 16182 19203 16216 19217
rect 16182 19183 16216 19203
rect 16278 19917 16312 19937
rect 16278 19903 16312 19917
rect 16278 19849 16312 19865
rect 16278 19831 16312 19849
rect 16278 19781 16312 19793
rect 16278 19759 16312 19781
rect 16278 19713 16312 19721
rect 16278 19687 16312 19713
rect 16278 19645 16312 19649
rect 16278 19615 16312 19645
rect 16278 19543 16312 19577
rect 16278 19475 16312 19505
rect 16278 19471 16312 19475
rect 16278 19407 16312 19433
rect 16278 19399 16312 19407
rect 16278 19339 16312 19361
rect 16278 19327 16312 19339
rect 16278 19271 16312 19289
rect 16278 19255 16312 19271
rect 16278 19203 16312 19217
rect 16278 19183 16312 19203
rect 16038 19088 16072 19122
rect 16230 19088 16264 19122
rect 13331 18836 13725 18942
rect 13900 18836 14294 18942
rect 16804 19265 16838 19299
rect 16804 19193 16838 19227
rect 16804 19121 16838 19155
rect 16804 19049 16838 19083
rect 16804 18977 16838 19011
rect 16804 18905 16838 18939
rect 17072 19198 17106 19232
rect 17144 19198 17178 19232
rect 13331 18450 13725 18556
rect 13900 18450 14294 18556
rect 13331 18064 13725 18170
rect 13900 18064 14294 18170
rect 15060 18532 15094 18566
rect 13331 17678 13725 17784
rect 13900 17678 14294 17784
rect 13331 17292 13725 17398
rect 13900 17292 14294 17398
rect 13331 16906 13725 17012
rect 13900 16906 14294 17012
rect 14660 17800 14694 17834
rect 14660 17728 14694 17762
rect 14660 17656 14694 17690
rect 14660 17584 14694 17618
rect 14660 17512 14694 17546
rect 14660 17440 14694 17474
rect 14660 17269 14694 17303
rect 14660 17197 14694 17231
rect 14660 17125 14694 17159
rect 14660 17053 14694 17087
rect 14660 16981 14694 17015
rect 14660 16909 14694 16943
rect 15016 18445 15050 18451
rect 15016 18417 15050 18445
rect 15016 18377 15050 18379
rect 15016 18345 15050 18377
rect 15016 18275 15050 18307
rect 15016 18273 15050 18275
rect 15016 18207 15050 18235
rect 15016 18201 15050 18207
rect 15016 18139 15050 18163
rect 15016 18129 15050 18139
rect 15016 18071 15050 18091
rect 15016 18057 15050 18071
rect 15016 18003 15050 18019
rect 15016 17985 15050 18003
rect 15016 17935 15050 17947
rect 15016 17913 15050 17935
rect 15016 17867 15050 17875
rect 15016 17841 15050 17867
rect 15016 17799 15050 17803
rect 15016 17769 15050 17799
rect 15016 17697 15050 17731
rect 15016 17629 15050 17659
rect 15016 17625 15050 17629
rect 15016 17561 15050 17587
rect 15016 17553 15050 17561
rect 15016 17493 15050 17515
rect 15016 17481 15050 17493
rect 15016 17425 15050 17443
rect 15016 17409 15050 17425
rect 15016 17357 15050 17371
rect 15016 17337 15050 17357
rect 15016 17289 15050 17299
rect 15016 17265 15050 17289
rect 15016 17221 15050 17227
rect 15016 17193 15050 17221
rect 15016 17153 15050 17155
rect 15016 17121 15050 17153
rect 15016 17051 15050 17083
rect 15016 17049 15050 17051
rect 15016 16983 15050 17011
rect 15016 16977 15050 16983
rect 15104 18445 15138 18451
rect 15104 18417 15138 18445
rect 15104 18377 15138 18379
rect 15104 18345 15138 18377
rect 15104 18275 15138 18307
rect 15104 18273 15138 18275
rect 15104 18207 15138 18235
rect 15104 18201 15138 18207
rect 15104 18139 15138 18163
rect 15104 18129 15138 18139
rect 15104 18071 15138 18091
rect 15104 18057 15138 18071
rect 15104 18003 15138 18019
rect 15104 17985 15138 18003
rect 15104 17935 15138 17947
rect 15104 17913 15138 17935
rect 15104 17867 15138 17875
rect 15104 17841 15138 17867
rect 15104 17799 15138 17803
rect 15104 17769 15138 17799
rect 15104 17697 15138 17731
rect 15104 17629 15138 17659
rect 15104 17625 15138 17629
rect 15104 17561 15138 17587
rect 15104 17553 15138 17561
rect 15104 17493 15138 17515
rect 15104 17481 15138 17493
rect 15104 17425 15138 17443
rect 15104 17409 15138 17425
rect 15104 17357 15138 17371
rect 15104 17337 15138 17357
rect 15104 17289 15138 17299
rect 15104 17265 15138 17289
rect 15104 17221 15138 17227
rect 15104 17193 15138 17221
rect 15104 17153 15138 17155
rect 15104 17121 15138 17153
rect 15104 17051 15138 17083
rect 15104 17049 15138 17051
rect 15104 16983 15138 17011
rect 15104 16977 15138 16983
rect 15470 18532 15504 18566
rect 15426 18445 15460 18451
rect 15426 18417 15460 18445
rect 15426 18377 15460 18379
rect 15426 18345 15460 18377
rect 15426 18275 15460 18307
rect 15426 18273 15460 18275
rect 15426 18207 15460 18235
rect 15426 18201 15460 18207
rect 15426 18139 15460 18163
rect 15426 18129 15460 18139
rect 15060 16862 15094 16896
rect 15426 18071 15460 18091
rect 15426 18057 15460 18071
rect 15426 18003 15460 18019
rect 15426 17985 15460 18003
rect 15426 17935 15460 17947
rect 15426 17913 15460 17935
rect 15426 17867 15460 17875
rect 15426 17841 15460 17867
rect 15426 17799 15460 17803
rect 15426 17769 15460 17799
rect 15426 17697 15460 17731
rect 15426 17629 15460 17659
rect 15426 17625 15460 17629
rect 15426 17561 15460 17587
rect 15426 17553 15460 17561
rect 15426 17493 15460 17515
rect 15426 17481 15460 17493
rect 15426 17425 15460 17443
rect 15426 17409 15460 17425
rect 15426 17357 15460 17371
rect 15426 17337 15460 17357
rect 15426 17289 15460 17299
rect 15426 17265 15460 17289
rect 15426 17221 15460 17227
rect 15426 17193 15460 17221
rect 15426 17153 15460 17155
rect 15426 17121 15460 17153
rect 15426 17051 15460 17083
rect 15426 17049 15460 17051
rect 15426 16983 15460 17011
rect 15426 16977 15460 16983
rect 15514 18445 15548 18451
rect 15514 18417 15548 18445
rect 15514 18377 15548 18379
rect 15514 18345 15548 18377
rect 15514 18275 15548 18307
rect 15514 18273 15548 18275
rect 15514 18207 15548 18235
rect 15514 18201 15548 18207
rect 15514 18139 15548 18163
rect 15514 18129 15548 18139
rect 15514 18071 15548 18091
rect 15514 18057 15548 18071
rect 15514 18003 15548 18019
rect 15514 17985 15548 18003
rect 15514 17935 15548 17947
rect 15514 17913 15548 17935
rect 15514 17867 15548 17875
rect 15514 17841 15548 17867
rect 15514 17799 15548 17803
rect 15514 17769 15548 17799
rect 15514 17697 15548 17731
rect 15514 17629 15548 17659
rect 15514 17625 15548 17629
rect 15514 17561 15548 17587
rect 15514 17553 15548 17561
rect 15514 17493 15548 17515
rect 15514 17481 15548 17493
rect 15514 17425 15548 17443
rect 15514 17409 15548 17425
rect 15514 17357 15548 17371
rect 15514 17337 15548 17357
rect 15514 17289 15548 17299
rect 15514 17265 15548 17289
rect 15514 17221 15548 17227
rect 15514 17193 15548 17221
rect 15514 17153 15548 17155
rect 15514 17121 15548 17153
rect 15514 17051 15548 17083
rect 15514 17049 15548 17051
rect 15514 16983 15548 17011
rect 15514 16977 15548 16983
rect 16272 18501 16306 18535
rect 16272 18429 16306 18463
rect 16272 18357 16306 18391
rect 16272 18285 16306 18319
rect 16272 18213 16306 18247
rect 16272 18141 16306 18175
rect 16816 18296 16850 18330
rect 15470 16862 15504 16896
rect 15880 17800 15914 17834
rect 15880 17728 15914 17762
rect 15880 17656 15914 17690
rect 15880 17584 15914 17618
rect 15880 17512 15914 17546
rect 15880 17440 15914 17474
rect 15880 17269 15914 17303
rect 15880 17197 15914 17231
rect 15880 17125 15914 17159
rect 15880 17053 15914 17087
rect 15880 16981 15914 17015
rect 15880 16909 15914 16943
rect 16272 17270 16306 17304
rect 16272 17198 16306 17232
rect 16272 17126 16306 17160
rect 16272 17054 16306 17088
rect 16272 16982 16306 17016
rect 16272 16910 16306 16944
rect 17414 21316 17448 21350
rect 17414 21244 17448 21278
rect 17414 21172 17448 21206
rect 17414 21100 17448 21134
rect 17414 21028 17448 21062
rect 17414 20956 17448 20990
rect 17414 17885 17448 17919
rect 17414 17813 17448 17847
rect 17414 17741 17448 17775
rect 17414 17669 17448 17703
rect 17414 17597 17448 17631
rect 17414 17525 17448 17559
rect 13338 16326 13444 16432
rect 14623 16367 14657 16401
rect 14695 16367 14729 16401
rect 15838 16367 15872 16401
rect 15910 16367 15944 16401
rect 14566 15942 14600 15976
rect 14758 15942 14792 15976
rect 14950 15942 14984 15976
rect 15142 15942 15176 15976
rect 13616 15502 13650 15536
rect 13572 15415 13606 15421
rect 13572 15387 13606 15415
rect 13572 15347 13606 15349
rect 13572 15315 13606 15347
rect 13660 15415 13694 15421
rect 13660 15387 13694 15415
rect 13660 15347 13694 15349
rect 13572 15245 13606 15277
rect 13572 15243 13606 15245
rect 13572 15177 13606 15205
rect 13572 15171 13606 15177
rect 13572 15109 13606 15133
rect 13572 15099 13606 15109
rect 13572 15041 13606 15061
rect 13572 15027 13606 15041
rect 13572 14973 13606 14989
rect 13572 14955 13606 14973
rect 13572 14905 13606 14917
rect 13572 14883 13606 14905
rect 13572 14837 13606 14845
rect 13572 14811 13606 14837
rect 13572 14769 13606 14773
rect 13572 14739 13606 14769
rect 13572 14667 13606 14701
rect 13572 14599 13606 14629
rect 13572 14595 13606 14599
rect 13572 14531 13606 14557
rect 13572 14523 13606 14531
rect 13572 14463 13606 14485
rect 13572 14451 13606 14463
rect 13572 14395 13606 14413
rect 13572 14379 13606 14395
rect 13572 14327 13606 14341
rect 13572 14307 13606 14327
rect 13572 14259 13606 14269
rect 13572 14235 13606 14259
rect 13572 14191 13606 14197
rect 13572 14163 13606 14191
rect 13572 14123 13606 14125
rect 13572 14091 13606 14123
rect 13572 14021 13606 14053
rect 13572 14019 13606 14021
rect 13572 13953 13606 13981
rect 13572 13947 13606 13953
rect 13660 15315 13694 15347
rect 13660 15245 13694 15277
rect 13660 15243 13694 15245
rect 13660 15177 13694 15205
rect 13660 15171 13694 15177
rect 13660 15109 13694 15133
rect 13660 15099 13694 15109
rect 13660 15041 13694 15061
rect 13660 15027 13694 15041
rect 13660 14973 13694 14989
rect 13660 14955 13694 14973
rect 13660 14905 13694 14917
rect 13660 14883 13694 14905
rect 13660 14837 13694 14845
rect 13660 14811 13694 14837
rect 13660 14769 13694 14773
rect 13660 14739 13694 14769
rect 13660 14667 13694 14701
rect 13660 14599 13694 14629
rect 13660 14595 13694 14599
rect 13660 14531 13694 14557
rect 13660 14523 13694 14531
rect 13660 14463 13694 14485
rect 13660 14451 13694 14463
rect 13660 14395 13694 14413
rect 13660 14379 13694 14395
rect 13660 14327 13694 14341
rect 13660 14307 13694 14327
rect 13660 14259 13694 14269
rect 13660 14235 13694 14259
rect 13660 14191 13694 14197
rect 13660 14163 13694 14191
rect 13660 14123 13694 14125
rect 13660 14091 13694 14123
rect 13660 14021 13694 14053
rect 13660 14019 13694 14021
rect 13660 13953 13694 13981
rect 13660 13947 13694 13953
rect 13616 13832 13650 13866
rect 14422 15839 14456 15857
rect 14422 15823 14456 15839
rect 14422 15771 14456 15785
rect 14422 15751 14456 15771
rect 14422 15703 14456 15713
rect 14422 15679 14456 15703
rect 14422 15635 14456 15641
rect 14422 15607 14456 15635
rect 14422 15567 14456 15569
rect 14422 15535 14456 15567
rect 14422 15465 14456 15497
rect 14422 15463 14456 15465
rect 14422 15397 14456 15425
rect 14422 15391 14456 15397
rect 14422 15329 14456 15353
rect 14422 15319 14456 15329
rect 14422 15261 14456 15281
rect 14422 15247 14456 15261
rect 14422 15193 14456 15209
rect 14422 15175 14456 15193
rect 14422 15125 14456 15137
rect 14422 15103 14456 15125
rect 14422 15057 14456 15065
rect 14422 15031 14456 15057
rect 14422 14989 14456 14993
rect 14422 14959 14456 14989
rect 14422 14887 14456 14921
rect 14422 14819 14456 14849
rect 14422 14815 14456 14819
rect 14422 14751 14456 14777
rect 14422 14743 14456 14751
rect 14422 14683 14456 14705
rect 14422 14671 14456 14683
rect 14422 14615 14456 14633
rect 14422 14599 14456 14615
rect 14422 14547 14456 14561
rect 14422 14527 14456 14547
rect 14422 14479 14456 14489
rect 14422 14455 14456 14479
rect 14422 14411 14456 14417
rect 14422 14383 14456 14411
rect 14422 14343 14456 14345
rect 14422 14311 14456 14343
rect 14422 14241 14456 14273
rect 14422 14239 14456 14241
rect 14422 14173 14456 14201
rect 14422 14167 14456 14173
rect 14422 14105 14456 14129
rect 14422 14095 14456 14105
rect 14422 14037 14456 14057
rect 14422 14023 14456 14037
rect 14422 13969 14456 13985
rect 14422 13951 14456 13969
rect 14518 15839 14552 15857
rect 14518 15823 14552 15839
rect 14518 15771 14552 15785
rect 14518 15751 14552 15771
rect 14518 15703 14552 15713
rect 14518 15679 14552 15703
rect 14518 15635 14552 15641
rect 14518 15607 14552 15635
rect 14518 15567 14552 15569
rect 14518 15535 14552 15567
rect 14518 15465 14552 15497
rect 14518 15463 14552 15465
rect 14518 15397 14552 15425
rect 14518 15391 14552 15397
rect 14518 15329 14552 15353
rect 14518 15319 14552 15329
rect 14518 15261 14552 15281
rect 14518 15247 14552 15261
rect 14518 15193 14552 15209
rect 14518 15175 14552 15193
rect 14518 15125 14552 15137
rect 14518 15103 14552 15125
rect 14518 15057 14552 15065
rect 14518 15031 14552 15057
rect 14518 14989 14552 14993
rect 14518 14959 14552 14989
rect 14518 14887 14552 14921
rect 14518 14819 14552 14849
rect 14518 14815 14552 14819
rect 14518 14751 14552 14777
rect 14518 14743 14552 14751
rect 14518 14683 14552 14705
rect 14518 14671 14552 14683
rect 14518 14615 14552 14633
rect 14518 14599 14552 14615
rect 14518 14547 14552 14561
rect 14518 14527 14552 14547
rect 14518 14479 14552 14489
rect 14518 14455 14552 14479
rect 14518 14411 14552 14417
rect 14518 14383 14552 14411
rect 14518 14343 14552 14345
rect 14518 14311 14552 14343
rect 14518 14241 14552 14273
rect 14518 14239 14552 14241
rect 14518 14173 14552 14201
rect 14518 14167 14552 14173
rect 14518 14105 14552 14129
rect 14518 14095 14552 14105
rect 14518 14037 14552 14057
rect 14518 14023 14552 14037
rect 14518 13969 14552 13985
rect 14518 13951 14552 13969
rect 14614 15839 14648 15857
rect 14614 15823 14648 15839
rect 14614 15771 14648 15785
rect 14614 15751 14648 15771
rect 14614 15703 14648 15713
rect 14614 15679 14648 15703
rect 14614 15635 14648 15641
rect 14614 15607 14648 15635
rect 14614 15567 14648 15569
rect 14614 15535 14648 15567
rect 14614 15465 14648 15497
rect 14614 15463 14648 15465
rect 14614 15397 14648 15425
rect 14614 15391 14648 15397
rect 14614 15329 14648 15353
rect 14614 15319 14648 15329
rect 14614 15261 14648 15281
rect 14614 15247 14648 15261
rect 14614 15193 14648 15209
rect 14614 15175 14648 15193
rect 14614 15125 14648 15137
rect 14614 15103 14648 15125
rect 14614 15057 14648 15065
rect 14614 15031 14648 15057
rect 14614 14989 14648 14993
rect 14614 14959 14648 14989
rect 14614 14887 14648 14921
rect 14614 14819 14648 14849
rect 14614 14815 14648 14819
rect 14614 14751 14648 14777
rect 14614 14743 14648 14751
rect 14614 14683 14648 14705
rect 14614 14671 14648 14683
rect 14614 14615 14648 14633
rect 14614 14599 14648 14615
rect 14614 14547 14648 14561
rect 14614 14527 14648 14547
rect 14614 14479 14648 14489
rect 14614 14455 14648 14479
rect 14614 14411 14648 14417
rect 14614 14383 14648 14411
rect 14614 14343 14648 14345
rect 14614 14311 14648 14343
rect 14614 14241 14648 14273
rect 14614 14239 14648 14241
rect 14614 14173 14648 14201
rect 14614 14167 14648 14173
rect 14614 14105 14648 14129
rect 14614 14095 14648 14105
rect 14614 14037 14648 14057
rect 14614 14023 14648 14037
rect 14614 13969 14648 13985
rect 14614 13951 14648 13969
rect 14710 15839 14744 15857
rect 14710 15823 14744 15839
rect 14710 15771 14744 15785
rect 14710 15751 14744 15771
rect 14710 15703 14744 15713
rect 14710 15679 14744 15703
rect 14710 15635 14744 15641
rect 14710 15607 14744 15635
rect 14710 15567 14744 15569
rect 14710 15535 14744 15567
rect 14710 15465 14744 15497
rect 14710 15463 14744 15465
rect 14710 15397 14744 15425
rect 14710 15391 14744 15397
rect 14710 15329 14744 15353
rect 14710 15319 14744 15329
rect 14710 15261 14744 15281
rect 14710 15247 14744 15261
rect 14710 15193 14744 15209
rect 14710 15175 14744 15193
rect 14710 15125 14744 15137
rect 14710 15103 14744 15125
rect 14710 15057 14744 15065
rect 14710 15031 14744 15057
rect 14710 14989 14744 14993
rect 14710 14959 14744 14989
rect 14710 14887 14744 14921
rect 14710 14819 14744 14849
rect 14710 14815 14744 14819
rect 14710 14751 14744 14777
rect 14710 14743 14744 14751
rect 14710 14683 14744 14705
rect 14710 14671 14744 14683
rect 14710 14615 14744 14633
rect 14710 14599 14744 14615
rect 14710 14547 14744 14561
rect 14710 14527 14744 14547
rect 14710 14479 14744 14489
rect 14710 14455 14744 14479
rect 14710 14411 14744 14417
rect 14710 14383 14744 14411
rect 14710 14343 14744 14345
rect 14710 14311 14744 14343
rect 14710 14241 14744 14273
rect 14710 14239 14744 14241
rect 14710 14173 14744 14201
rect 14710 14167 14744 14173
rect 14710 14105 14744 14129
rect 14710 14095 14744 14105
rect 14710 14037 14744 14057
rect 14710 14023 14744 14037
rect 14710 13969 14744 13985
rect 14710 13951 14744 13969
rect 14806 15839 14840 15857
rect 14806 15823 14840 15839
rect 14806 15771 14840 15785
rect 14806 15751 14840 15771
rect 14806 15703 14840 15713
rect 14806 15679 14840 15703
rect 14806 15635 14840 15641
rect 14806 15607 14840 15635
rect 14806 15567 14840 15569
rect 14806 15535 14840 15567
rect 14806 15465 14840 15497
rect 14806 15463 14840 15465
rect 14806 15397 14840 15425
rect 14806 15391 14840 15397
rect 14806 15329 14840 15353
rect 14806 15319 14840 15329
rect 14806 15261 14840 15281
rect 14806 15247 14840 15261
rect 14806 15193 14840 15209
rect 14806 15175 14840 15193
rect 14806 15125 14840 15137
rect 14806 15103 14840 15125
rect 14806 15057 14840 15065
rect 14806 15031 14840 15057
rect 14806 14989 14840 14993
rect 14806 14959 14840 14989
rect 14806 14887 14840 14921
rect 14806 14819 14840 14849
rect 14806 14815 14840 14819
rect 14806 14751 14840 14777
rect 14806 14743 14840 14751
rect 14806 14683 14840 14705
rect 14806 14671 14840 14683
rect 14806 14615 14840 14633
rect 14806 14599 14840 14615
rect 14806 14547 14840 14561
rect 14806 14527 14840 14547
rect 14806 14479 14840 14489
rect 14806 14455 14840 14479
rect 14806 14411 14840 14417
rect 14806 14383 14840 14411
rect 14806 14343 14840 14345
rect 14806 14311 14840 14343
rect 14806 14241 14840 14273
rect 14806 14239 14840 14241
rect 14806 14173 14840 14201
rect 14806 14167 14840 14173
rect 14806 14105 14840 14129
rect 14806 14095 14840 14105
rect 14806 14037 14840 14057
rect 14806 14023 14840 14037
rect 14806 13969 14840 13985
rect 14806 13951 14840 13969
rect 14902 15839 14936 15857
rect 14902 15823 14936 15839
rect 14902 15771 14936 15785
rect 14902 15751 14936 15771
rect 14902 15703 14936 15713
rect 14902 15679 14936 15703
rect 14902 15635 14936 15641
rect 14902 15607 14936 15635
rect 14902 15567 14936 15569
rect 14902 15535 14936 15567
rect 14902 15465 14936 15497
rect 14902 15463 14936 15465
rect 14902 15397 14936 15425
rect 14902 15391 14936 15397
rect 14902 15329 14936 15353
rect 14902 15319 14936 15329
rect 14902 15261 14936 15281
rect 14902 15247 14936 15261
rect 14902 15193 14936 15209
rect 14902 15175 14936 15193
rect 14902 15125 14936 15137
rect 14902 15103 14936 15125
rect 14902 15057 14936 15065
rect 14902 15031 14936 15057
rect 14902 14989 14936 14993
rect 14902 14959 14936 14989
rect 14902 14887 14936 14921
rect 14902 14819 14936 14849
rect 14902 14815 14936 14819
rect 14902 14751 14936 14777
rect 14902 14743 14936 14751
rect 14902 14683 14936 14705
rect 14902 14671 14936 14683
rect 14902 14615 14936 14633
rect 14902 14599 14936 14615
rect 14902 14547 14936 14561
rect 14902 14527 14936 14547
rect 14902 14479 14936 14489
rect 14902 14455 14936 14479
rect 14902 14411 14936 14417
rect 14902 14383 14936 14411
rect 14902 14343 14936 14345
rect 14902 14311 14936 14343
rect 14902 14241 14936 14273
rect 14902 14239 14936 14241
rect 14902 14173 14936 14201
rect 14902 14167 14936 14173
rect 14902 14105 14936 14129
rect 14902 14095 14936 14105
rect 14902 14037 14936 14057
rect 14902 14023 14936 14037
rect 14902 13969 14936 13985
rect 14902 13951 14936 13969
rect 14998 15839 15032 15857
rect 14998 15823 15032 15839
rect 14998 15771 15032 15785
rect 14998 15751 15032 15771
rect 14998 15703 15032 15713
rect 14998 15679 15032 15703
rect 14998 15635 15032 15641
rect 14998 15607 15032 15635
rect 14998 15567 15032 15569
rect 14998 15535 15032 15567
rect 14998 15465 15032 15497
rect 14998 15463 15032 15465
rect 14998 15397 15032 15425
rect 14998 15391 15032 15397
rect 14998 15329 15032 15353
rect 14998 15319 15032 15329
rect 14998 15261 15032 15281
rect 14998 15247 15032 15261
rect 14998 15193 15032 15209
rect 14998 15175 15032 15193
rect 14998 15125 15032 15137
rect 14998 15103 15032 15125
rect 14998 15057 15032 15065
rect 14998 15031 15032 15057
rect 14998 14989 15032 14993
rect 14998 14959 15032 14989
rect 14998 14887 15032 14921
rect 14998 14819 15032 14849
rect 14998 14815 15032 14819
rect 14998 14751 15032 14777
rect 14998 14743 15032 14751
rect 14998 14683 15032 14705
rect 14998 14671 15032 14683
rect 14998 14615 15032 14633
rect 14998 14599 15032 14615
rect 14998 14547 15032 14561
rect 14998 14527 15032 14547
rect 14998 14479 15032 14489
rect 14998 14455 15032 14479
rect 14998 14411 15032 14417
rect 14998 14383 15032 14411
rect 14998 14343 15032 14345
rect 14998 14311 15032 14343
rect 14998 14241 15032 14273
rect 14998 14239 15032 14241
rect 14998 14173 15032 14201
rect 14998 14167 15032 14173
rect 14998 14105 15032 14129
rect 14998 14095 15032 14105
rect 14998 14037 15032 14057
rect 14998 14023 15032 14037
rect 14998 13969 15032 13985
rect 14998 13951 15032 13969
rect 15094 15839 15128 15857
rect 15094 15823 15128 15839
rect 15094 15771 15128 15785
rect 15094 15751 15128 15771
rect 15094 15703 15128 15713
rect 15094 15679 15128 15703
rect 15094 15635 15128 15641
rect 15094 15607 15128 15635
rect 15094 15567 15128 15569
rect 15094 15535 15128 15567
rect 15094 15465 15128 15497
rect 15094 15463 15128 15465
rect 15094 15397 15128 15425
rect 15094 15391 15128 15397
rect 15094 15329 15128 15353
rect 15094 15319 15128 15329
rect 15094 15261 15128 15281
rect 15094 15247 15128 15261
rect 15094 15193 15128 15209
rect 15094 15175 15128 15193
rect 15094 15125 15128 15137
rect 15094 15103 15128 15125
rect 15094 15057 15128 15065
rect 15094 15031 15128 15057
rect 15094 14989 15128 14993
rect 15094 14959 15128 14989
rect 15094 14887 15128 14921
rect 15094 14819 15128 14849
rect 15094 14815 15128 14819
rect 15094 14751 15128 14777
rect 15094 14743 15128 14751
rect 15094 14683 15128 14705
rect 15094 14671 15128 14683
rect 15094 14615 15128 14633
rect 15094 14599 15128 14615
rect 15094 14547 15128 14561
rect 15094 14527 15128 14547
rect 15094 14479 15128 14489
rect 15094 14455 15128 14479
rect 15094 14411 15128 14417
rect 15094 14383 15128 14411
rect 15094 14343 15128 14345
rect 15094 14311 15128 14343
rect 15094 14241 15128 14273
rect 15094 14239 15128 14241
rect 15094 14173 15128 14201
rect 15094 14167 15128 14173
rect 15094 14105 15128 14129
rect 15094 14095 15128 14105
rect 15094 14037 15128 14057
rect 15094 14023 15128 14037
rect 15094 13969 15128 13985
rect 15094 13951 15128 13969
rect 15190 15839 15224 15857
rect 15190 15823 15224 15839
rect 15190 15771 15224 15785
rect 15190 15751 15224 15771
rect 15190 15703 15224 15713
rect 15190 15679 15224 15703
rect 15190 15635 15224 15641
rect 15190 15607 15224 15635
rect 15190 15567 15224 15569
rect 15190 15535 15224 15567
rect 15190 15465 15224 15497
rect 15190 15463 15224 15465
rect 15190 15397 15224 15425
rect 15190 15391 15224 15397
rect 15190 15329 15224 15353
rect 15190 15319 15224 15329
rect 15190 15261 15224 15281
rect 15190 15247 15224 15261
rect 15190 15193 15224 15209
rect 15190 15175 15224 15193
rect 15190 15125 15224 15137
rect 15190 15103 15224 15125
rect 15190 15057 15224 15065
rect 15190 15031 15224 15057
rect 15190 14989 15224 14993
rect 15190 14959 15224 14989
rect 15190 14887 15224 14921
rect 15190 14819 15224 14849
rect 15190 14815 15224 14819
rect 15190 14751 15224 14777
rect 15190 14743 15224 14751
rect 15190 14683 15224 14705
rect 15190 14671 15224 14683
rect 15190 14615 15224 14633
rect 15190 14599 15224 14615
rect 15190 14547 15224 14561
rect 15190 14527 15224 14547
rect 15190 14479 15224 14489
rect 15190 14455 15224 14479
rect 15190 14411 15224 14417
rect 15190 14383 15224 14411
rect 15190 14343 15224 14345
rect 15190 14311 15224 14343
rect 15190 14241 15224 14273
rect 15190 14239 15224 14241
rect 15190 14173 15224 14201
rect 15190 14167 15224 14173
rect 15190 14105 15224 14129
rect 15190 14095 15224 14105
rect 15190 14037 15224 14057
rect 15190 14023 15224 14037
rect 15190 13969 15224 13985
rect 15190 13951 15224 13969
rect 14470 13832 14504 13866
rect 14662 13832 14696 13866
rect 14854 13832 14888 13866
rect 15046 13832 15080 13866
rect 16166 15910 16200 15944
rect 16166 15838 16200 15872
rect 16166 15766 16200 15800
rect 16166 15694 16200 15728
rect 16166 15622 16200 15656
rect 16166 15550 16200 15584
rect 16166 14239 16200 14273
rect 16166 14167 16200 14201
rect 16166 14095 16200 14129
rect 16166 14023 16200 14057
rect 16166 13951 16200 13985
rect 16166 13879 16200 13913
rect 17236 15990 17270 16024
rect 17092 15878 17126 15896
rect 17092 15862 17126 15878
rect 17092 15810 17126 15824
rect 17092 15790 17126 15810
rect 17092 15742 17126 15752
rect 17092 15718 17126 15742
rect 17092 15674 17126 15680
rect 17092 15646 17126 15674
rect 17092 15606 17126 15608
rect 17092 15574 17126 15606
rect 17092 15504 17126 15536
rect 17092 15502 17126 15504
rect 17092 15436 17126 15464
rect 17092 15430 17126 15436
rect 17092 15368 17126 15392
rect 17092 15358 17126 15368
rect 17092 15300 17126 15320
rect 17092 15286 17126 15300
rect 17092 15232 17126 15248
rect 17092 15214 17126 15232
rect 17092 15164 17126 15176
rect 17092 15142 17126 15164
rect 17092 15096 17126 15104
rect 17092 15070 17126 15096
rect 17092 15028 17126 15032
rect 17092 14998 17126 15028
rect 17092 14926 17126 14960
rect 17092 14858 17126 14888
rect 17092 14854 17126 14858
rect 17092 14790 17126 14816
rect 17092 14782 17126 14790
rect 17092 14722 17126 14744
rect 17092 14710 17126 14722
rect 17092 14654 17126 14672
rect 17092 14638 17126 14654
rect 17092 14586 17126 14600
rect 17092 14566 17126 14586
rect 17092 14518 17126 14528
rect 17092 14494 17126 14518
rect 17092 14450 17126 14456
rect 17092 14422 17126 14450
rect 17092 14382 17126 14384
rect 17092 14350 17126 14382
rect 17092 14280 17126 14312
rect 17092 14278 17126 14280
rect 17092 14212 17126 14240
rect 17092 14206 17126 14212
rect 17092 14144 17126 14168
rect 17092 14134 17126 14144
rect 17092 14076 17126 14096
rect 17092 14062 17126 14076
rect 17092 14008 17126 14024
rect 17092 13990 17126 14008
rect 17188 15878 17222 15896
rect 17188 15862 17222 15878
rect 17188 15810 17222 15824
rect 17188 15790 17222 15810
rect 17188 15742 17222 15752
rect 17188 15718 17222 15742
rect 17188 15674 17222 15680
rect 17188 15646 17222 15674
rect 17188 15606 17222 15608
rect 17188 15574 17222 15606
rect 17188 15504 17222 15536
rect 17188 15502 17222 15504
rect 17188 15436 17222 15464
rect 17188 15430 17222 15436
rect 17188 15368 17222 15392
rect 17188 15358 17222 15368
rect 17188 15300 17222 15320
rect 17188 15286 17222 15300
rect 17188 15232 17222 15248
rect 17188 15214 17222 15232
rect 17188 15164 17222 15176
rect 17188 15142 17222 15164
rect 17188 15096 17222 15104
rect 17188 15070 17222 15096
rect 17188 15028 17222 15032
rect 17188 14998 17222 15028
rect 17188 14926 17222 14960
rect 17188 14858 17222 14888
rect 17188 14854 17222 14858
rect 17188 14790 17222 14816
rect 17188 14782 17222 14790
rect 17188 14722 17222 14744
rect 17188 14710 17222 14722
rect 17188 14654 17222 14672
rect 17188 14638 17222 14654
rect 17188 14586 17222 14600
rect 17188 14566 17222 14586
rect 17188 14518 17222 14528
rect 17188 14494 17222 14518
rect 17188 14450 17222 14456
rect 17188 14422 17222 14450
rect 17188 14382 17222 14384
rect 17188 14350 17222 14382
rect 17188 14280 17222 14312
rect 17188 14278 17222 14280
rect 17188 14212 17222 14240
rect 17188 14206 17222 14212
rect 17188 14144 17222 14168
rect 17188 14134 17222 14144
rect 17188 14076 17222 14096
rect 17188 14062 17222 14076
rect 17188 14008 17222 14024
rect 17188 13990 17222 14008
rect 17284 15878 17318 15896
rect 17284 15862 17318 15878
rect 17380 15878 17414 15896
rect 17380 15862 17414 15878
rect 17284 15810 17318 15824
rect 17284 15790 17318 15810
rect 17284 15742 17318 15752
rect 17284 15718 17318 15742
rect 17284 15674 17318 15680
rect 17284 15646 17318 15674
rect 17284 15606 17318 15608
rect 17284 15574 17318 15606
rect 17284 15504 17318 15536
rect 17284 15502 17318 15504
rect 17284 15436 17318 15464
rect 17284 15430 17318 15436
rect 17284 15368 17318 15392
rect 17284 15358 17318 15368
rect 17284 15300 17318 15320
rect 17284 15286 17318 15300
rect 17284 15232 17318 15248
rect 17284 15214 17318 15232
rect 17284 15164 17318 15176
rect 17284 15142 17318 15164
rect 17284 15096 17318 15104
rect 17284 15070 17318 15096
rect 17284 15028 17318 15032
rect 17284 14998 17318 15028
rect 17284 14926 17318 14960
rect 17284 14858 17318 14888
rect 17284 14854 17318 14858
rect 17284 14790 17318 14816
rect 17284 14782 17318 14790
rect 17284 14722 17318 14744
rect 17284 14710 17318 14722
rect 17284 14654 17318 14672
rect 17284 14638 17318 14654
rect 17284 14586 17318 14600
rect 17284 14566 17318 14586
rect 17284 14518 17318 14528
rect 17284 14494 17318 14518
rect 17284 14450 17318 14456
rect 17284 14422 17318 14450
rect 17284 14382 17318 14384
rect 17284 14350 17318 14382
rect 17284 14280 17318 14312
rect 17284 14278 17318 14280
rect 17284 14212 17318 14240
rect 17284 14206 17318 14212
rect 17284 14144 17318 14168
rect 17284 14134 17318 14144
rect 17284 14076 17318 14096
rect 17284 14062 17318 14076
rect 17284 14008 17318 14024
rect 17284 13990 17318 14008
rect 17380 15810 17414 15824
rect 17380 15790 17414 15810
rect 17380 15742 17414 15752
rect 17380 15718 17414 15742
rect 17380 15674 17414 15680
rect 17380 15646 17414 15674
rect 17380 15606 17414 15608
rect 17380 15574 17414 15606
rect 17380 15504 17414 15536
rect 17380 15502 17414 15504
rect 17380 15436 17414 15464
rect 17380 15430 17414 15436
rect 17380 15368 17414 15392
rect 17380 15358 17414 15368
rect 17380 15300 17414 15320
rect 17380 15286 17414 15300
rect 17380 15232 17414 15248
rect 17380 15214 17414 15232
rect 17380 15164 17414 15176
rect 17380 15142 17414 15164
rect 17380 15096 17414 15104
rect 17380 15070 17414 15096
rect 17380 15028 17414 15032
rect 17380 14998 17414 15028
rect 17380 14926 17414 14960
rect 17380 14858 17414 14888
rect 17380 14854 17414 14858
rect 17380 14790 17414 14816
rect 17380 14782 17414 14790
rect 17380 14722 17414 14744
rect 17380 14710 17414 14722
rect 17380 14654 17414 14672
rect 17380 14638 17414 14654
rect 17380 14586 17414 14600
rect 17380 14566 17414 14586
rect 17380 14518 17414 14528
rect 17380 14494 17414 14518
rect 17380 14450 17414 14456
rect 17380 14422 17414 14450
rect 17380 14382 17414 14384
rect 17380 14350 17414 14382
rect 17380 14280 17414 14312
rect 17380 14278 17414 14280
rect 17380 14212 17414 14240
rect 17380 14206 17414 14212
rect 17380 14144 17414 14168
rect 17380 14134 17414 14144
rect 17380 14076 17414 14096
rect 17380 14062 17414 14076
rect 17380 14008 17414 14024
rect 17380 13990 17414 14008
rect 17140 13862 17174 13896
rect 17332 13862 17366 13896
rect 16165 13297 16199 13331
rect 17040 13276 17074 13310
rect 13509 13147 13543 13181
rect 13434 13005 13468 13023
rect 13434 12989 13468 13005
rect 13434 12937 13468 12951
rect 13434 12917 13468 12937
rect 13434 12869 13468 12879
rect 13434 12845 13468 12869
rect 13434 12801 13468 12807
rect 13434 12773 13468 12801
rect 13434 12733 13468 12735
rect 13434 12701 13468 12733
rect 13434 12631 13468 12663
rect 13434 12629 13468 12631
rect 13434 12563 13468 12591
rect 13434 12557 13468 12563
rect 13434 12495 13468 12519
rect 13434 12485 13468 12495
rect 13434 12427 13468 12447
rect 13434 12413 13468 12427
rect 13434 12359 13468 12375
rect 13434 12341 13468 12359
rect 13434 12291 13468 12303
rect 13434 12269 13468 12291
rect 13434 12223 13468 12231
rect 13434 12197 13468 12223
rect 13434 12155 13468 12159
rect 13434 12125 13468 12155
rect 13434 12053 13468 12087
rect 13434 11985 13468 12015
rect 13434 11981 13468 11985
rect 13434 11917 13468 11943
rect 13434 11909 13468 11917
rect 13434 11849 13468 11871
rect 13434 11837 13468 11849
rect 13434 11781 13468 11799
rect 13434 11765 13468 11781
rect 13434 11713 13468 11727
rect 13434 11693 13468 11713
rect 13434 11645 13468 11655
rect 13434 11621 13468 11645
rect 13434 11577 13468 11583
rect 13434 11549 13468 11577
rect 13434 11509 13468 11511
rect 13434 11477 13468 11509
rect 13434 11407 13468 11439
rect 13434 11405 13468 11407
rect 13434 11339 13468 11367
rect 13434 11333 13468 11339
rect 13434 11271 13468 11295
rect 13434 11261 13468 11271
rect 13434 11203 13468 11223
rect 13434 11189 13468 11203
rect 13434 11135 13468 11151
rect 13434 11117 13468 11135
rect 13522 13005 13556 13023
rect 13522 12989 13556 13005
rect 13522 12937 13556 12951
rect 13522 12917 13556 12937
rect 13522 12869 13556 12879
rect 13522 12845 13556 12869
rect 13522 12801 13556 12807
rect 13522 12773 13556 12801
rect 13522 12733 13556 12735
rect 13522 12701 13556 12733
rect 13522 12631 13556 12663
rect 13522 12629 13556 12631
rect 13522 12563 13556 12591
rect 13522 12557 13556 12563
rect 13522 12495 13556 12519
rect 13522 12485 13556 12495
rect 13522 12427 13556 12447
rect 13522 12413 13556 12427
rect 13522 12359 13556 12375
rect 13522 12341 13556 12359
rect 13522 12291 13556 12303
rect 13522 12269 13556 12291
rect 13522 12223 13556 12231
rect 13522 12197 13556 12223
rect 13522 12155 13556 12159
rect 13522 12125 13556 12155
rect 13522 12053 13556 12087
rect 13522 11985 13556 12015
rect 13522 11981 13556 11985
rect 13522 11917 13556 11943
rect 13522 11909 13556 11917
rect 13522 11849 13556 11871
rect 13522 11837 13556 11849
rect 13522 11781 13556 11799
rect 13522 11765 13556 11781
rect 13522 11713 13556 11727
rect 13522 11693 13556 11713
rect 13522 11645 13556 11655
rect 13522 11621 13556 11645
rect 13522 11577 13556 11583
rect 13522 11549 13556 11577
rect 13522 11509 13556 11511
rect 13522 11477 13556 11509
rect 13522 11407 13556 11439
rect 13522 11405 13556 11407
rect 13522 11339 13556 11367
rect 13522 11333 13556 11339
rect 13522 11271 13556 11295
rect 13522 11261 13556 11271
rect 13522 11203 13556 11223
rect 13522 11189 13556 11203
rect 13522 11135 13556 11151
rect 13522 11117 13556 11135
rect 13610 13005 13644 13023
rect 13610 12989 13644 13005
rect 13610 12937 13644 12951
rect 13610 12917 13644 12937
rect 13610 12869 13644 12879
rect 13610 12845 13644 12869
rect 13610 12801 13644 12807
rect 13610 12773 13644 12801
rect 13610 12733 13644 12735
rect 13610 12701 13644 12733
rect 13610 12631 13644 12663
rect 13610 12629 13644 12631
rect 13610 12563 13644 12591
rect 13610 12557 13644 12563
rect 13610 12495 13644 12519
rect 13610 12485 13644 12495
rect 13610 12427 13644 12447
rect 13610 12413 13644 12427
rect 13610 12359 13644 12375
rect 13610 12341 13644 12359
rect 13610 12291 13644 12303
rect 13610 12269 13644 12291
rect 13610 12223 13644 12231
rect 13610 12197 13644 12223
rect 13610 12155 13644 12159
rect 13610 12125 13644 12155
rect 13610 12053 13644 12087
rect 13610 11985 13644 12015
rect 13610 11981 13644 11985
rect 13610 11917 13644 11943
rect 13610 11909 13644 11917
rect 13610 11849 13644 11871
rect 13610 11837 13644 11849
rect 13610 11781 13644 11799
rect 13610 11765 13644 11781
rect 13610 11713 13644 11727
rect 13610 11693 13644 11713
rect 13610 11645 13644 11655
rect 13610 11621 13644 11645
rect 13610 11577 13644 11583
rect 13610 11549 13644 11577
rect 13610 11509 13644 11511
rect 13610 11477 13644 11509
rect 13610 11407 13644 11439
rect 13610 11405 13644 11407
rect 13610 11339 13644 11367
rect 13610 11333 13644 11339
rect 13610 11271 13644 11295
rect 13610 11261 13644 11271
rect 13610 11203 13644 11223
rect 13610 11189 13644 11203
rect 13610 11135 13644 11151
rect 13610 11117 13644 11135
rect 13698 13005 13732 13023
rect 13698 12989 13732 13005
rect 13698 12937 13732 12951
rect 13698 12917 13732 12937
rect 13698 12869 13732 12879
rect 13698 12845 13732 12869
rect 13698 12801 13732 12807
rect 13698 12773 13732 12801
rect 13698 12733 13732 12735
rect 13698 12701 13732 12733
rect 13698 12631 13732 12663
rect 13698 12629 13732 12631
rect 13698 12563 13732 12591
rect 13698 12557 13732 12563
rect 13698 12495 13732 12519
rect 13698 12485 13732 12495
rect 13698 12427 13732 12447
rect 13698 12413 13732 12427
rect 13698 12359 13732 12375
rect 13698 12341 13732 12359
rect 13698 12291 13732 12303
rect 13698 12269 13732 12291
rect 13698 12223 13732 12231
rect 13698 12197 13732 12223
rect 13698 12155 13732 12159
rect 13698 12125 13732 12155
rect 13698 12053 13732 12087
rect 13698 11985 13732 12015
rect 13698 11981 13732 11985
rect 13698 11917 13732 11943
rect 13698 11909 13732 11917
rect 13698 11849 13732 11871
rect 13698 11837 13732 11849
rect 13698 11781 13732 11799
rect 13698 11765 13732 11781
rect 13698 11713 13732 11727
rect 13698 11693 13732 11713
rect 13698 11645 13732 11655
rect 13698 11621 13732 11645
rect 13698 11577 13732 11583
rect 13698 11549 13732 11577
rect 13698 11509 13732 11511
rect 13698 11477 13732 11509
rect 13698 11407 13732 11439
rect 13698 11405 13732 11407
rect 13698 11339 13732 11367
rect 13698 11333 13732 11339
rect 13698 11271 13732 11295
rect 13698 11261 13732 11271
rect 13698 11203 13732 11223
rect 13698 11189 13732 11203
rect 13698 11135 13732 11151
rect 13698 11117 13732 11135
rect 13786 13005 13820 13023
rect 13786 12989 13820 13005
rect 13786 12937 13820 12951
rect 13786 12917 13820 12937
rect 13786 12869 13820 12879
rect 13786 12845 13820 12869
rect 13786 12801 13820 12807
rect 13786 12773 13820 12801
rect 13786 12733 13820 12735
rect 13786 12701 13820 12733
rect 13786 12631 13820 12663
rect 13786 12629 13820 12631
rect 13786 12563 13820 12591
rect 13786 12557 13820 12563
rect 13786 12495 13820 12519
rect 13786 12485 13820 12495
rect 13786 12427 13820 12447
rect 13786 12413 13820 12427
rect 13786 12359 13820 12375
rect 13786 12341 13820 12359
rect 13786 12291 13820 12303
rect 13786 12269 13820 12291
rect 13786 12223 13820 12231
rect 13786 12197 13820 12223
rect 13786 12155 13820 12159
rect 13786 12125 13820 12155
rect 13786 12053 13820 12087
rect 13786 11985 13820 12015
rect 13786 11981 13820 11985
rect 13786 11917 13820 11943
rect 13786 11909 13820 11917
rect 13786 11849 13820 11871
rect 13786 11837 13820 11849
rect 13786 11781 13820 11799
rect 13786 11765 13820 11781
rect 13786 11713 13820 11727
rect 13786 11693 13820 11713
rect 13786 11645 13820 11655
rect 13786 11621 13820 11645
rect 13786 11577 13820 11583
rect 13786 11549 13820 11577
rect 13786 11509 13820 11511
rect 13786 11477 13820 11509
rect 13786 11407 13820 11439
rect 13786 11405 13820 11407
rect 13786 11339 13820 11367
rect 13786 11333 13820 11339
rect 13786 11271 13820 11295
rect 13786 11261 13820 11271
rect 13786 11203 13820 11223
rect 13786 11189 13820 11203
rect 13786 11135 13820 11151
rect 13786 11117 13820 11135
rect 13874 13005 13908 13023
rect 13874 12989 13908 13005
rect 13874 12937 13908 12951
rect 13874 12917 13908 12937
rect 13874 12869 13908 12879
rect 13874 12845 13908 12869
rect 13874 12801 13908 12807
rect 13874 12773 13908 12801
rect 13874 12733 13908 12735
rect 13874 12701 13908 12733
rect 13874 12631 13908 12663
rect 13874 12629 13908 12631
rect 13874 12563 13908 12591
rect 13874 12557 13908 12563
rect 13874 12495 13908 12519
rect 13874 12485 13908 12495
rect 13874 12427 13908 12447
rect 13874 12413 13908 12427
rect 13874 12359 13908 12375
rect 13874 12341 13908 12359
rect 13874 12291 13908 12303
rect 13874 12269 13908 12291
rect 13874 12223 13908 12231
rect 13874 12197 13908 12223
rect 13874 12155 13908 12159
rect 13874 12125 13908 12155
rect 13874 12053 13908 12087
rect 13874 11985 13908 12015
rect 13874 11981 13908 11985
rect 13874 11917 13908 11943
rect 13874 11909 13908 11917
rect 13874 11849 13908 11871
rect 13874 11837 13908 11849
rect 13874 11781 13908 11799
rect 13874 11765 13908 11781
rect 13874 11713 13908 11727
rect 13874 11693 13908 11713
rect 13874 11645 13908 11655
rect 13874 11621 13908 11645
rect 13874 11577 13908 11583
rect 13874 11549 13908 11577
rect 13874 11509 13908 11511
rect 13874 11477 13908 11509
rect 13874 11407 13908 11439
rect 13874 11405 13908 11407
rect 13874 11339 13908 11367
rect 13874 11333 13908 11339
rect 13874 11271 13908 11295
rect 13874 11261 13908 11271
rect 13874 11203 13908 11223
rect 13874 11189 13908 11203
rect 13874 11135 13908 11151
rect 13874 11117 13908 11135
rect 13962 13005 13996 13023
rect 13962 12989 13996 13005
rect 13962 12937 13996 12951
rect 13962 12917 13996 12937
rect 13962 12869 13996 12879
rect 13962 12845 13996 12869
rect 13962 12801 13996 12807
rect 13962 12773 13996 12801
rect 13962 12733 13996 12735
rect 13962 12701 13996 12733
rect 13962 12631 13996 12663
rect 13962 12629 13996 12631
rect 13962 12563 13996 12591
rect 13962 12557 13996 12563
rect 13962 12495 13996 12519
rect 13962 12485 13996 12495
rect 13962 12427 13996 12447
rect 13962 12413 13996 12427
rect 13962 12359 13996 12375
rect 13962 12341 13996 12359
rect 13962 12291 13996 12303
rect 13962 12269 13996 12291
rect 13962 12223 13996 12231
rect 13962 12197 13996 12223
rect 13962 12155 13996 12159
rect 13962 12125 13996 12155
rect 13962 12053 13996 12087
rect 13962 11985 13996 12015
rect 13962 11981 13996 11985
rect 13962 11917 13996 11943
rect 13962 11909 13996 11917
rect 13962 11849 13996 11871
rect 13962 11837 13996 11849
rect 13962 11781 13996 11799
rect 13962 11765 13996 11781
rect 13962 11713 13996 11727
rect 13962 11693 13996 11713
rect 13962 11645 13996 11655
rect 13962 11621 13996 11645
rect 13962 11577 13996 11583
rect 13962 11549 13996 11577
rect 13962 11509 13996 11511
rect 13962 11477 13996 11509
rect 13962 11407 13996 11439
rect 13962 11405 13996 11407
rect 13962 11339 13996 11367
rect 13962 11333 13996 11339
rect 13962 11271 13996 11295
rect 13962 11261 13996 11271
rect 13962 11203 13996 11223
rect 13962 11189 13996 11203
rect 13962 11135 13996 11151
rect 13962 11117 13996 11135
rect 14050 13005 14084 13023
rect 14050 12989 14084 13005
rect 14050 12937 14084 12951
rect 14050 12917 14084 12937
rect 14050 12869 14084 12879
rect 14050 12845 14084 12869
rect 14050 12801 14084 12807
rect 14050 12773 14084 12801
rect 14050 12733 14084 12735
rect 14050 12701 14084 12733
rect 14050 12631 14084 12663
rect 14050 12629 14084 12631
rect 14050 12563 14084 12591
rect 14050 12557 14084 12563
rect 14050 12495 14084 12519
rect 14050 12485 14084 12495
rect 14050 12427 14084 12447
rect 14050 12413 14084 12427
rect 14050 12359 14084 12375
rect 14050 12341 14084 12359
rect 14050 12291 14084 12303
rect 14050 12269 14084 12291
rect 14050 12223 14084 12231
rect 14050 12197 14084 12223
rect 14050 12155 14084 12159
rect 14050 12125 14084 12155
rect 14050 12053 14084 12087
rect 14050 11985 14084 12015
rect 14050 11981 14084 11985
rect 14050 11917 14084 11943
rect 14050 11909 14084 11917
rect 14050 11849 14084 11871
rect 14050 11837 14084 11849
rect 14050 11781 14084 11799
rect 14050 11765 14084 11781
rect 14050 11713 14084 11727
rect 14050 11693 14084 11713
rect 14050 11645 14084 11655
rect 14050 11621 14084 11645
rect 14050 11577 14084 11583
rect 14050 11549 14084 11577
rect 14050 11509 14084 11511
rect 14050 11477 14084 11509
rect 14050 11407 14084 11439
rect 14050 11405 14084 11407
rect 14050 11339 14084 11367
rect 14050 11333 14084 11339
rect 14050 11271 14084 11295
rect 14050 11261 14084 11271
rect 14050 11203 14084 11223
rect 14050 11189 14084 11203
rect 14050 11135 14084 11151
rect 14050 11117 14084 11135
rect 14138 13005 14172 13023
rect 14138 12989 14172 13005
rect 14138 12937 14172 12951
rect 14138 12917 14172 12937
rect 14138 12869 14172 12879
rect 14138 12845 14172 12869
rect 14138 12801 14172 12807
rect 14138 12773 14172 12801
rect 14138 12733 14172 12735
rect 14138 12701 14172 12733
rect 14138 12631 14172 12663
rect 14138 12629 14172 12631
rect 14138 12563 14172 12591
rect 14138 12557 14172 12563
rect 14138 12495 14172 12519
rect 14138 12485 14172 12495
rect 14138 12427 14172 12447
rect 14138 12413 14172 12427
rect 14138 12359 14172 12375
rect 14138 12341 14172 12359
rect 14138 12291 14172 12303
rect 14138 12269 14172 12291
rect 14138 12223 14172 12231
rect 14138 12197 14172 12223
rect 14138 12155 14172 12159
rect 14138 12125 14172 12155
rect 14138 12053 14172 12087
rect 14138 11985 14172 12015
rect 14138 11981 14172 11985
rect 14138 11917 14172 11943
rect 14138 11909 14172 11917
rect 14138 11849 14172 11871
rect 14138 11837 14172 11849
rect 14138 11781 14172 11799
rect 14138 11765 14172 11781
rect 14138 11713 14172 11727
rect 14138 11693 14172 11713
rect 14138 11645 14172 11655
rect 14138 11621 14172 11645
rect 14138 11577 14172 11583
rect 14138 11549 14172 11577
rect 14138 11509 14172 11511
rect 14138 11477 14172 11509
rect 14138 11407 14172 11439
rect 14138 11405 14172 11407
rect 14138 11339 14172 11367
rect 14138 11333 14172 11339
rect 14138 11271 14172 11295
rect 14138 11261 14172 11271
rect 14138 11203 14172 11223
rect 14138 11189 14172 11203
rect 14138 11135 14172 11151
rect 14138 11117 14172 11135
rect 14226 13005 14260 13023
rect 14226 12989 14260 13005
rect 14226 12937 14260 12951
rect 14226 12917 14260 12937
rect 14226 12869 14260 12879
rect 14226 12845 14260 12869
rect 14226 12801 14260 12807
rect 14226 12773 14260 12801
rect 14226 12733 14260 12735
rect 14226 12701 14260 12733
rect 14226 12631 14260 12663
rect 14226 12629 14260 12631
rect 14226 12563 14260 12591
rect 14226 12557 14260 12563
rect 14226 12495 14260 12519
rect 14226 12485 14260 12495
rect 14226 12427 14260 12447
rect 14226 12413 14260 12427
rect 14226 12359 14260 12375
rect 14226 12341 14260 12359
rect 14226 12291 14260 12303
rect 14226 12269 14260 12291
rect 14226 12223 14260 12231
rect 14226 12197 14260 12223
rect 14226 12155 14260 12159
rect 14226 12125 14260 12155
rect 14226 12053 14260 12087
rect 14226 11985 14260 12015
rect 14226 11981 14260 11985
rect 14226 11917 14260 11943
rect 14226 11909 14260 11917
rect 14226 11849 14260 11871
rect 14226 11837 14260 11849
rect 14226 11781 14260 11799
rect 14226 11765 14260 11781
rect 14226 11713 14260 11727
rect 14226 11693 14260 11713
rect 14226 11645 14260 11655
rect 14226 11621 14260 11645
rect 14226 11577 14260 11583
rect 14226 11549 14260 11577
rect 14226 11509 14260 11511
rect 14226 11477 14260 11509
rect 14226 11407 14260 11439
rect 14226 11405 14260 11407
rect 14226 11339 14260 11367
rect 14226 11333 14260 11339
rect 14226 11271 14260 11295
rect 14226 11261 14260 11271
rect 14226 11203 14260 11223
rect 14226 11189 14260 11203
rect 14226 11135 14260 11151
rect 14226 11117 14260 11135
rect 14314 13005 14348 13023
rect 14314 12989 14348 13005
rect 14314 12937 14348 12951
rect 14314 12917 14348 12937
rect 14314 12869 14348 12879
rect 14314 12845 14348 12869
rect 14314 12801 14348 12807
rect 14314 12773 14348 12801
rect 14314 12733 14348 12735
rect 14314 12701 14348 12733
rect 14314 12631 14348 12663
rect 14314 12629 14348 12631
rect 14314 12563 14348 12591
rect 14314 12557 14348 12563
rect 14314 12495 14348 12519
rect 14314 12485 14348 12495
rect 14314 12427 14348 12447
rect 14314 12413 14348 12427
rect 14314 12359 14348 12375
rect 14314 12341 14348 12359
rect 14314 12291 14348 12303
rect 14314 12269 14348 12291
rect 14314 12223 14348 12231
rect 14314 12197 14348 12223
rect 14314 12155 14348 12159
rect 14314 12125 14348 12155
rect 14314 12053 14348 12087
rect 14314 11985 14348 12015
rect 14314 11981 14348 11985
rect 14314 11917 14348 11943
rect 14314 11909 14348 11917
rect 14314 11849 14348 11871
rect 14314 11837 14348 11849
rect 14314 11781 14348 11799
rect 14314 11765 14348 11781
rect 14314 11713 14348 11727
rect 14314 11693 14348 11713
rect 14314 11645 14348 11655
rect 14314 11621 14348 11645
rect 14314 11577 14348 11583
rect 14314 11549 14348 11577
rect 14314 11509 14348 11511
rect 14314 11477 14348 11509
rect 14314 11407 14348 11439
rect 14314 11405 14348 11407
rect 14314 11339 14348 11367
rect 14314 11333 14348 11339
rect 14314 11271 14348 11295
rect 14314 11261 14348 11271
rect 14314 11203 14348 11223
rect 14314 11189 14348 11203
rect 14314 11135 14348 11151
rect 14314 11117 14348 11135
rect 14402 13005 14436 13023
rect 14402 12989 14436 13005
rect 14402 12937 14436 12951
rect 14402 12917 14436 12937
rect 14402 12869 14436 12879
rect 14402 12845 14436 12869
rect 14402 12801 14436 12807
rect 14402 12773 14436 12801
rect 14402 12733 14436 12735
rect 14402 12701 14436 12733
rect 14402 12631 14436 12663
rect 14402 12629 14436 12631
rect 14402 12563 14436 12591
rect 14402 12557 14436 12563
rect 14402 12495 14436 12519
rect 14402 12485 14436 12495
rect 14402 12427 14436 12447
rect 14402 12413 14436 12427
rect 14402 12359 14436 12375
rect 14402 12341 14436 12359
rect 14402 12291 14436 12303
rect 14402 12269 14436 12291
rect 14402 12223 14436 12231
rect 14402 12197 14436 12223
rect 14402 12155 14436 12159
rect 14402 12125 14436 12155
rect 14402 12053 14436 12087
rect 14402 11985 14436 12015
rect 14402 11981 14436 11985
rect 14402 11917 14436 11943
rect 14402 11909 14436 11917
rect 14402 11849 14436 11871
rect 14402 11837 14436 11849
rect 14402 11781 14436 11799
rect 14402 11765 14436 11781
rect 14402 11713 14436 11727
rect 14402 11693 14436 11713
rect 14402 11645 14436 11655
rect 14402 11621 14436 11645
rect 14402 11577 14436 11583
rect 14402 11549 14436 11577
rect 14402 11509 14436 11511
rect 14402 11477 14436 11509
rect 14402 11407 14436 11439
rect 14402 11405 14436 11407
rect 14402 11339 14436 11367
rect 14402 11333 14436 11339
rect 14402 11271 14436 11295
rect 14402 11261 14436 11271
rect 14402 11203 14436 11223
rect 14402 11189 14436 11203
rect 14402 11135 14436 11151
rect 14402 11117 14436 11135
rect 14490 13005 14524 13023
rect 14490 12989 14524 13005
rect 14490 12937 14524 12951
rect 14490 12917 14524 12937
rect 14490 12869 14524 12879
rect 14490 12845 14524 12869
rect 14490 12801 14524 12807
rect 14490 12773 14524 12801
rect 14490 12733 14524 12735
rect 14490 12701 14524 12733
rect 14490 12631 14524 12663
rect 14490 12629 14524 12631
rect 14490 12563 14524 12591
rect 14490 12557 14524 12563
rect 14490 12495 14524 12519
rect 14490 12485 14524 12495
rect 14490 12427 14524 12447
rect 14490 12413 14524 12427
rect 14490 12359 14524 12375
rect 14490 12341 14524 12359
rect 14490 12291 14524 12303
rect 14490 12269 14524 12291
rect 14490 12223 14524 12231
rect 14490 12197 14524 12223
rect 14490 12155 14524 12159
rect 14490 12125 14524 12155
rect 14490 12053 14524 12087
rect 14490 11985 14524 12015
rect 14490 11981 14524 11985
rect 14490 11917 14524 11943
rect 14490 11909 14524 11917
rect 14490 11849 14524 11871
rect 14490 11837 14524 11849
rect 14490 11781 14524 11799
rect 14490 11765 14524 11781
rect 14490 11713 14524 11727
rect 14490 11693 14524 11713
rect 14490 11645 14524 11655
rect 14490 11621 14524 11645
rect 14490 11577 14524 11583
rect 14490 11549 14524 11577
rect 14490 11509 14524 11511
rect 14490 11477 14524 11509
rect 14490 11407 14524 11439
rect 14490 11405 14524 11407
rect 14490 11339 14524 11367
rect 14490 11333 14524 11339
rect 14490 11271 14524 11295
rect 14490 11261 14524 11271
rect 14490 11203 14524 11223
rect 14490 11189 14524 11203
rect 14490 11135 14524 11151
rect 14490 11117 14524 11135
rect 14578 13005 14612 13023
rect 14578 12989 14612 13005
rect 14578 12937 14612 12951
rect 14578 12917 14612 12937
rect 14578 12869 14612 12879
rect 14578 12845 14612 12869
rect 14578 12801 14612 12807
rect 14578 12773 14612 12801
rect 14578 12733 14612 12735
rect 14578 12701 14612 12733
rect 14578 12631 14612 12663
rect 14578 12629 14612 12631
rect 14578 12563 14612 12591
rect 14578 12557 14612 12563
rect 14578 12495 14612 12519
rect 14578 12485 14612 12495
rect 14578 12427 14612 12447
rect 14578 12413 14612 12427
rect 14578 12359 14612 12375
rect 14578 12341 14612 12359
rect 14578 12291 14612 12303
rect 14578 12269 14612 12291
rect 14578 12223 14612 12231
rect 14578 12197 14612 12223
rect 14578 12155 14612 12159
rect 14578 12125 14612 12155
rect 14578 12053 14612 12087
rect 14578 11985 14612 12015
rect 14578 11981 14612 11985
rect 14578 11917 14612 11943
rect 14578 11909 14612 11917
rect 14578 11849 14612 11871
rect 14578 11837 14612 11849
rect 14578 11781 14612 11799
rect 14578 11765 14612 11781
rect 14578 11713 14612 11727
rect 14578 11693 14612 11713
rect 14578 11645 14612 11655
rect 14578 11621 14612 11645
rect 14578 11577 14612 11583
rect 14578 11549 14612 11577
rect 14578 11509 14612 11511
rect 14578 11477 14612 11509
rect 14578 11407 14612 11439
rect 14578 11405 14612 11407
rect 14578 11339 14612 11367
rect 14578 11333 14612 11339
rect 14578 11271 14612 11295
rect 14578 11261 14612 11271
rect 14578 11203 14612 11223
rect 14578 11189 14612 11203
rect 14578 11135 14612 11151
rect 14578 11117 14612 11135
rect 14666 13005 14700 13023
rect 14666 12989 14700 13005
rect 14666 12937 14700 12951
rect 14666 12917 14700 12937
rect 14666 12869 14700 12879
rect 14666 12845 14700 12869
rect 14666 12801 14700 12807
rect 14666 12773 14700 12801
rect 14666 12733 14700 12735
rect 14666 12701 14700 12733
rect 14666 12631 14700 12663
rect 14666 12629 14700 12631
rect 14666 12563 14700 12591
rect 14666 12557 14700 12563
rect 14666 12495 14700 12519
rect 14666 12485 14700 12495
rect 14666 12427 14700 12447
rect 14666 12413 14700 12427
rect 14666 12359 14700 12375
rect 14666 12341 14700 12359
rect 14666 12291 14700 12303
rect 14666 12269 14700 12291
rect 14666 12223 14700 12231
rect 14666 12197 14700 12223
rect 14666 12155 14700 12159
rect 14666 12125 14700 12155
rect 14666 12053 14700 12087
rect 14666 11985 14700 12015
rect 14666 11981 14700 11985
rect 14666 11917 14700 11943
rect 14666 11909 14700 11917
rect 14666 11849 14700 11871
rect 14666 11837 14700 11849
rect 14666 11781 14700 11799
rect 14666 11765 14700 11781
rect 14666 11713 14700 11727
rect 14666 11693 14700 11713
rect 14666 11645 14700 11655
rect 14666 11621 14700 11645
rect 14666 11577 14700 11583
rect 14666 11549 14700 11577
rect 14666 11509 14700 11511
rect 14666 11477 14700 11509
rect 14666 11407 14700 11439
rect 14666 11405 14700 11407
rect 14666 11339 14700 11367
rect 14666 11333 14700 11339
rect 14666 11271 14700 11295
rect 14666 11261 14700 11271
rect 14666 11203 14700 11223
rect 14666 11189 14700 11203
rect 14666 11135 14700 11151
rect 14666 11117 14700 11135
rect 14754 13005 14788 13023
rect 14754 12989 14788 13005
rect 14754 12937 14788 12951
rect 14754 12917 14788 12937
rect 14754 12869 14788 12879
rect 14754 12845 14788 12869
rect 14754 12801 14788 12807
rect 14754 12773 14788 12801
rect 14754 12733 14788 12735
rect 14754 12701 14788 12733
rect 14754 12631 14788 12663
rect 14754 12629 14788 12631
rect 14754 12563 14788 12591
rect 14754 12557 14788 12563
rect 14754 12495 14788 12519
rect 14754 12485 14788 12495
rect 14754 12427 14788 12447
rect 14754 12413 14788 12427
rect 14754 12359 14788 12375
rect 14754 12341 14788 12359
rect 14754 12291 14788 12303
rect 14754 12269 14788 12291
rect 14754 12223 14788 12231
rect 14754 12197 14788 12223
rect 14754 12155 14788 12159
rect 14754 12125 14788 12155
rect 14754 12053 14788 12087
rect 14754 11985 14788 12015
rect 14754 11981 14788 11985
rect 14754 11917 14788 11943
rect 14754 11909 14788 11917
rect 14754 11849 14788 11871
rect 14754 11837 14788 11849
rect 14754 11781 14788 11799
rect 14754 11765 14788 11781
rect 14754 11713 14788 11727
rect 14754 11693 14788 11713
rect 14754 11645 14788 11655
rect 14754 11621 14788 11645
rect 14754 11577 14788 11583
rect 14754 11549 14788 11577
rect 14754 11509 14788 11511
rect 14754 11477 14788 11509
rect 14754 11407 14788 11439
rect 14754 11405 14788 11407
rect 14754 11339 14788 11367
rect 14754 11333 14788 11339
rect 14754 11271 14788 11295
rect 14754 11261 14788 11271
rect 14754 11203 14788 11223
rect 14754 11189 14788 11203
rect 14754 11135 14788 11151
rect 14754 11117 14788 11135
rect 14842 13005 14876 13023
rect 14842 12989 14876 13005
rect 14842 12937 14876 12951
rect 14842 12917 14876 12937
rect 14842 12869 14876 12879
rect 14842 12845 14876 12869
rect 14842 12801 14876 12807
rect 14842 12773 14876 12801
rect 14842 12733 14876 12735
rect 14842 12701 14876 12733
rect 14842 12631 14876 12663
rect 14842 12629 14876 12631
rect 14842 12563 14876 12591
rect 14842 12557 14876 12563
rect 14842 12495 14876 12519
rect 14842 12485 14876 12495
rect 14842 12427 14876 12447
rect 14842 12413 14876 12427
rect 14842 12359 14876 12375
rect 14842 12341 14876 12359
rect 14842 12291 14876 12303
rect 14842 12269 14876 12291
rect 14842 12223 14876 12231
rect 14842 12197 14876 12223
rect 14842 12155 14876 12159
rect 14842 12125 14876 12155
rect 14842 12053 14876 12087
rect 14842 11985 14876 12015
rect 14842 11981 14876 11985
rect 14842 11917 14876 11943
rect 14842 11909 14876 11917
rect 14842 11849 14876 11871
rect 14842 11837 14876 11849
rect 14842 11781 14876 11799
rect 14842 11765 14876 11781
rect 14842 11713 14876 11727
rect 14842 11693 14876 11713
rect 14842 11645 14876 11655
rect 14842 11621 14876 11645
rect 14842 11577 14876 11583
rect 14842 11549 14876 11577
rect 14842 11509 14876 11511
rect 14842 11477 14876 11509
rect 14842 11407 14876 11439
rect 14842 11405 14876 11407
rect 14842 11339 14876 11367
rect 14842 11333 14876 11339
rect 14842 11271 14876 11295
rect 14842 11261 14876 11271
rect 14842 11203 14876 11223
rect 14842 11189 14876 11203
rect 14842 11135 14876 11151
rect 14842 11117 14876 11135
rect 14930 13005 14964 13023
rect 14930 12989 14964 13005
rect 14930 12937 14964 12951
rect 14930 12917 14964 12937
rect 14930 12869 14964 12879
rect 14930 12845 14964 12869
rect 14930 12801 14964 12807
rect 14930 12773 14964 12801
rect 14930 12733 14964 12735
rect 14930 12701 14964 12733
rect 14930 12631 14964 12663
rect 14930 12629 14964 12631
rect 14930 12563 14964 12591
rect 14930 12557 14964 12563
rect 14930 12495 14964 12519
rect 14930 12485 14964 12495
rect 14930 12427 14964 12447
rect 14930 12413 14964 12427
rect 14930 12359 14964 12375
rect 14930 12341 14964 12359
rect 14930 12291 14964 12303
rect 14930 12269 14964 12291
rect 14930 12223 14964 12231
rect 14930 12197 14964 12223
rect 14930 12155 14964 12159
rect 14930 12125 14964 12155
rect 14930 12053 14964 12087
rect 14930 11985 14964 12015
rect 14930 11981 14964 11985
rect 14930 11917 14964 11943
rect 14930 11909 14964 11917
rect 14930 11849 14964 11871
rect 14930 11837 14964 11849
rect 14930 11781 14964 11799
rect 14930 11765 14964 11781
rect 14930 11713 14964 11727
rect 14930 11693 14964 11713
rect 14930 11645 14964 11655
rect 14930 11621 14964 11645
rect 14930 11577 14964 11583
rect 14930 11549 14964 11577
rect 14930 11509 14964 11511
rect 14930 11477 14964 11509
rect 14930 11407 14964 11439
rect 14930 11405 14964 11407
rect 14930 11339 14964 11367
rect 14930 11333 14964 11339
rect 14930 11271 14964 11295
rect 14930 11261 14964 11271
rect 14930 11203 14964 11223
rect 14930 11189 14964 11203
rect 14930 11135 14964 11151
rect 14930 11117 14964 11135
rect 15018 13005 15052 13023
rect 15018 12989 15052 13005
rect 15018 12937 15052 12951
rect 15018 12917 15052 12937
rect 15018 12869 15052 12879
rect 15018 12845 15052 12869
rect 15018 12801 15052 12807
rect 15018 12773 15052 12801
rect 15018 12733 15052 12735
rect 15018 12701 15052 12733
rect 15018 12631 15052 12663
rect 15018 12629 15052 12631
rect 15018 12563 15052 12591
rect 15018 12557 15052 12563
rect 15018 12495 15052 12519
rect 15018 12485 15052 12495
rect 15018 12427 15052 12447
rect 15018 12413 15052 12427
rect 15018 12359 15052 12375
rect 15018 12341 15052 12359
rect 15018 12291 15052 12303
rect 15018 12269 15052 12291
rect 15018 12223 15052 12231
rect 15018 12197 15052 12223
rect 15018 12155 15052 12159
rect 15018 12125 15052 12155
rect 15018 12053 15052 12087
rect 15018 11985 15052 12015
rect 15018 11981 15052 11985
rect 15018 11917 15052 11943
rect 15018 11909 15052 11917
rect 15018 11849 15052 11871
rect 15018 11837 15052 11849
rect 15018 11781 15052 11799
rect 15018 11765 15052 11781
rect 15018 11713 15052 11727
rect 15018 11693 15052 11713
rect 15018 11645 15052 11655
rect 15018 11621 15052 11645
rect 15018 11577 15052 11583
rect 15018 11549 15052 11577
rect 15018 11509 15052 11511
rect 15018 11477 15052 11509
rect 15018 11407 15052 11439
rect 15018 11405 15052 11407
rect 15018 11339 15052 11367
rect 15018 11333 15052 11339
rect 15018 11271 15052 11295
rect 15018 11261 15052 11271
rect 15018 11203 15052 11223
rect 15018 11189 15052 11203
rect 15018 11135 15052 11151
rect 15018 11117 15052 11135
rect 15106 13005 15140 13023
rect 15106 12989 15140 13005
rect 15106 12937 15140 12951
rect 15106 12917 15140 12937
rect 15106 12869 15140 12879
rect 15106 12845 15140 12869
rect 15106 12801 15140 12807
rect 15106 12773 15140 12801
rect 15106 12733 15140 12735
rect 15106 12701 15140 12733
rect 15106 12631 15140 12663
rect 15106 12629 15140 12631
rect 15106 12563 15140 12591
rect 15106 12557 15140 12563
rect 15106 12495 15140 12519
rect 15106 12485 15140 12495
rect 15106 12427 15140 12447
rect 15106 12413 15140 12427
rect 15106 12359 15140 12375
rect 15106 12341 15140 12359
rect 15106 12291 15140 12303
rect 15106 12269 15140 12291
rect 15106 12223 15140 12231
rect 15106 12197 15140 12223
rect 15106 12155 15140 12159
rect 15106 12125 15140 12155
rect 15106 12053 15140 12087
rect 15106 11985 15140 12015
rect 15106 11981 15140 11985
rect 15106 11917 15140 11943
rect 15106 11909 15140 11917
rect 15106 11849 15140 11871
rect 15106 11837 15140 11849
rect 15106 11781 15140 11799
rect 15106 11765 15140 11781
rect 15106 11713 15140 11727
rect 15106 11693 15140 11713
rect 15106 11645 15140 11655
rect 15106 11621 15140 11645
rect 15106 11577 15140 11583
rect 15106 11549 15140 11577
rect 15106 11509 15140 11511
rect 15106 11477 15140 11509
rect 15106 11407 15140 11439
rect 15106 11405 15140 11407
rect 15106 11339 15140 11367
rect 15106 11333 15140 11339
rect 15106 11271 15140 11295
rect 15106 11261 15140 11271
rect 15106 11203 15140 11223
rect 15106 11189 15140 11203
rect 15106 11135 15140 11151
rect 15106 11117 15140 11135
rect 15194 13005 15228 13023
rect 15194 12989 15228 13005
rect 15194 12937 15228 12951
rect 15194 12917 15228 12937
rect 15194 12869 15228 12879
rect 15194 12845 15228 12869
rect 15194 12801 15228 12807
rect 15194 12773 15228 12801
rect 15194 12733 15228 12735
rect 15194 12701 15228 12733
rect 15194 12631 15228 12663
rect 15194 12629 15228 12631
rect 15194 12563 15228 12591
rect 15194 12557 15228 12563
rect 15194 12495 15228 12519
rect 15194 12485 15228 12495
rect 15194 12427 15228 12447
rect 15194 12413 15228 12427
rect 15194 12359 15228 12375
rect 15194 12341 15228 12359
rect 15194 12291 15228 12303
rect 15194 12269 15228 12291
rect 15194 12223 15228 12231
rect 15194 12197 15228 12223
rect 15194 12155 15228 12159
rect 15194 12125 15228 12155
rect 15194 12053 15228 12087
rect 15194 11985 15228 12015
rect 15194 11981 15228 11985
rect 15194 11917 15228 11943
rect 15194 11909 15228 11917
rect 15194 11849 15228 11871
rect 15194 11837 15228 11849
rect 15194 11781 15228 11799
rect 15194 11765 15228 11781
rect 15194 11713 15228 11727
rect 15194 11693 15228 11713
rect 15194 11645 15228 11655
rect 15194 11621 15228 11645
rect 15194 11577 15228 11583
rect 15194 11549 15228 11577
rect 15194 11509 15228 11511
rect 15194 11477 15228 11509
rect 15194 11407 15228 11439
rect 15194 11405 15228 11407
rect 15194 11339 15228 11367
rect 15194 11333 15228 11339
rect 15194 11271 15228 11295
rect 15194 11261 15228 11271
rect 15194 11203 15228 11223
rect 15194 11189 15228 11203
rect 15194 11135 15228 11151
rect 15194 11117 15228 11135
rect 15282 13005 15316 13023
rect 15282 12989 15316 13005
rect 15282 12937 15316 12951
rect 15282 12917 15316 12937
rect 15282 12869 15316 12879
rect 15282 12845 15316 12869
rect 15282 12801 15316 12807
rect 15282 12773 15316 12801
rect 15282 12733 15316 12735
rect 15282 12701 15316 12733
rect 15282 12631 15316 12663
rect 15282 12629 15316 12631
rect 15282 12563 15316 12591
rect 15282 12557 15316 12563
rect 15282 12495 15316 12519
rect 15282 12485 15316 12495
rect 15282 12427 15316 12447
rect 15282 12413 15316 12427
rect 15282 12359 15316 12375
rect 15282 12341 15316 12359
rect 15282 12291 15316 12303
rect 15282 12269 15316 12291
rect 15282 12223 15316 12231
rect 15282 12197 15316 12223
rect 15282 12155 15316 12159
rect 15282 12125 15316 12155
rect 15282 12053 15316 12087
rect 15282 11985 15316 12015
rect 15282 11981 15316 11985
rect 15282 11917 15316 11943
rect 15282 11909 15316 11917
rect 15282 11849 15316 11871
rect 15282 11837 15316 11849
rect 15282 11781 15316 11799
rect 15282 11765 15316 11781
rect 15282 11713 15316 11727
rect 15282 11693 15316 11713
rect 15282 11645 15316 11655
rect 15282 11621 15316 11645
rect 15282 11577 15316 11583
rect 15282 11549 15316 11577
rect 15282 11509 15316 11511
rect 15282 11477 15316 11509
rect 15282 11407 15316 11439
rect 15282 11405 15316 11407
rect 15282 11339 15316 11367
rect 15282 11333 15316 11339
rect 15282 11271 15316 11295
rect 15282 11261 15316 11271
rect 15282 11203 15316 11223
rect 15282 11189 15316 11203
rect 15282 11135 15316 11151
rect 15282 11117 15316 11135
rect 15370 13005 15404 13023
rect 15370 12989 15404 13005
rect 15370 12937 15404 12951
rect 15370 12917 15404 12937
rect 15370 12869 15404 12879
rect 15370 12845 15404 12869
rect 15370 12801 15404 12807
rect 15370 12773 15404 12801
rect 15370 12733 15404 12735
rect 15370 12701 15404 12733
rect 15370 12631 15404 12663
rect 15370 12629 15404 12631
rect 15370 12563 15404 12591
rect 15370 12557 15404 12563
rect 15370 12495 15404 12519
rect 15370 12485 15404 12495
rect 15370 12427 15404 12447
rect 15370 12413 15404 12427
rect 15370 12359 15404 12375
rect 15370 12341 15404 12359
rect 15370 12291 15404 12303
rect 15370 12269 15404 12291
rect 15370 12223 15404 12231
rect 15370 12197 15404 12223
rect 15370 12155 15404 12159
rect 15370 12125 15404 12155
rect 15370 12053 15404 12087
rect 15370 11985 15404 12015
rect 15370 11981 15404 11985
rect 15370 11917 15404 11943
rect 15370 11909 15404 11917
rect 15370 11849 15404 11871
rect 15370 11837 15404 11849
rect 15370 11781 15404 11799
rect 15370 11765 15404 11781
rect 15370 11713 15404 11727
rect 15370 11693 15404 11713
rect 15370 11645 15404 11655
rect 15370 11621 15404 11645
rect 15370 11577 15404 11583
rect 15370 11549 15404 11577
rect 15370 11509 15404 11511
rect 15370 11477 15404 11509
rect 15370 11407 15404 11439
rect 15370 11405 15404 11407
rect 15370 11339 15404 11367
rect 15370 11333 15404 11339
rect 15370 11271 15404 11295
rect 15370 11261 15404 11271
rect 15370 11203 15404 11223
rect 15370 11189 15404 11203
rect 15370 11135 15404 11151
rect 15370 11117 15404 11135
rect 15458 13005 15492 13023
rect 15458 12989 15492 13005
rect 15458 12937 15492 12951
rect 15458 12917 15492 12937
rect 15458 12869 15492 12879
rect 15458 12845 15492 12869
rect 15458 12801 15492 12807
rect 15458 12773 15492 12801
rect 15458 12733 15492 12735
rect 15458 12701 15492 12733
rect 15458 12631 15492 12663
rect 15458 12629 15492 12631
rect 15458 12563 15492 12591
rect 15458 12557 15492 12563
rect 15458 12495 15492 12519
rect 15458 12485 15492 12495
rect 15458 12427 15492 12447
rect 15458 12413 15492 12427
rect 15458 12359 15492 12375
rect 15458 12341 15492 12359
rect 15458 12291 15492 12303
rect 15458 12269 15492 12291
rect 15458 12223 15492 12231
rect 15458 12197 15492 12223
rect 15458 12155 15492 12159
rect 15458 12125 15492 12155
rect 15458 12053 15492 12087
rect 15458 11985 15492 12015
rect 15458 11981 15492 11985
rect 15458 11917 15492 11943
rect 15458 11909 15492 11917
rect 15458 11849 15492 11871
rect 15458 11837 15492 11849
rect 15458 11781 15492 11799
rect 15458 11765 15492 11781
rect 15458 11713 15492 11727
rect 15458 11693 15492 11713
rect 15458 11645 15492 11655
rect 15458 11621 15492 11645
rect 15458 11577 15492 11583
rect 15458 11549 15492 11577
rect 15458 11509 15492 11511
rect 15458 11477 15492 11509
rect 15458 11407 15492 11439
rect 15458 11405 15492 11407
rect 15458 11339 15492 11367
rect 15458 11333 15492 11339
rect 15458 11271 15492 11295
rect 15458 11261 15492 11271
rect 15458 11203 15492 11223
rect 15458 11189 15492 11203
rect 15458 11135 15492 11151
rect 15458 11117 15492 11135
rect 15546 13005 15580 13023
rect 15546 12989 15580 13005
rect 15546 12937 15580 12951
rect 15546 12917 15580 12937
rect 15546 12869 15580 12879
rect 15546 12845 15580 12869
rect 15546 12801 15580 12807
rect 15546 12773 15580 12801
rect 15546 12733 15580 12735
rect 15546 12701 15580 12733
rect 15546 12631 15580 12663
rect 15546 12629 15580 12631
rect 15546 12563 15580 12591
rect 15546 12557 15580 12563
rect 15546 12495 15580 12519
rect 15546 12485 15580 12495
rect 15546 12427 15580 12447
rect 15546 12413 15580 12427
rect 15546 12359 15580 12375
rect 15546 12341 15580 12359
rect 15546 12291 15580 12303
rect 15546 12269 15580 12291
rect 15546 12223 15580 12231
rect 15546 12197 15580 12223
rect 15546 12155 15580 12159
rect 15546 12125 15580 12155
rect 15546 12053 15580 12087
rect 15546 11985 15580 12015
rect 15546 11981 15580 11985
rect 15546 11917 15580 11943
rect 15546 11909 15580 11917
rect 15546 11849 15580 11871
rect 15546 11837 15580 11849
rect 15546 11781 15580 11799
rect 15546 11765 15580 11781
rect 15546 11713 15580 11727
rect 15546 11693 15580 11713
rect 15546 11645 15580 11655
rect 15546 11621 15580 11645
rect 15546 11577 15580 11583
rect 15546 11549 15580 11577
rect 15546 11509 15580 11511
rect 15546 11477 15580 11509
rect 15546 11407 15580 11439
rect 15546 11405 15580 11407
rect 15546 11339 15580 11367
rect 15546 11333 15580 11339
rect 15546 11271 15580 11295
rect 15546 11261 15580 11271
rect 15546 11203 15580 11223
rect 15546 11189 15580 11203
rect 15546 11135 15580 11151
rect 15546 11117 15580 11135
rect 15634 13005 15668 13023
rect 15634 12989 15668 13005
rect 15634 12937 15668 12951
rect 15634 12917 15668 12937
rect 15634 12869 15668 12879
rect 15634 12845 15668 12869
rect 15634 12801 15668 12807
rect 15634 12773 15668 12801
rect 15634 12733 15668 12735
rect 15634 12701 15668 12733
rect 15634 12631 15668 12663
rect 15634 12629 15668 12631
rect 15634 12563 15668 12591
rect 15634 12557 15668 12563
rect 15634 12495 15668 12519
rect 15634 12485 15668 12495
rect 15634 12427 15668 12447
rect 15634 12413 15668 12427
rect 15634 12359 15668 12375
rect 15634 12341 15668 12359
rect 15634 12291 15668 12303
rect 15634 12269 15668 12291
rect 15634 12223 15668 12231
rect 15634 12197 15668 12223
rect 15634 12155 15668 12159
rect 15634 12125 15668 12155
rect 15634 12053 15668 12087
rect 15634 11985 15668 12015
rect 15634 11981 15668 11985
rect 15634 11917 15668 11943
rect 15634 11909 15668 11917
rect 15634 11849 15668 11871
rect 15634 11837 15668 11849
rect 15634 11781 15668 11799
rect 15634 11765 15668 11781
rect 15634 11713 15668 11727
rect 15634 11693 15668 11713
rect 15634 11645 15668 11655
rect 15634 11621 15668 11645
rect 15634 11577 15668 11583
rect 15634 11549 15668 11577
rect 15634 11509 15668 11511
rect 15634 11477 15668 11509
rect 15634 11407 15668 11439
rect 15634 11405 15668 11407
rect 15634 11339 15668 11367
rect 15634 11333 15668 11339
rect 15634 11271 15668 11295
rect 15634 11261 15668 11271
rect 15634 11203 15668 11223
rect 15634 11189 15668 11203
rect 15634 11135 15668 11151
rect 15634 11117 15668 11135
rect 15722 13005 15756 13023
rect 15722 12989 15756 13005
rect 15722 12937 15756 12951
rect 15722 12917 15756 12937
rect 15722 12869 15756 12879
rect 15722 12845 15756 12869
rect 15722 12801 15756 12807
rect 15722 12773 15756 12801
rect 15722 12733 15756 12735
rect 15722 12701 15756 12733
rect 15722 12631 15756 12663
rect 15722 12629 15756 12631
rect 15722 12563 15756 12591
rect 15722 12557 15756 12563
rect 15722 12495 15756 12519
rect 15722 12485 15756 12495
rect 15722 12427 15756 12447
rect 15722 12413 15756 12427
rect 15722 12359 15756 12375
rect 15722 12341 15756 12359
rect 15722 12291 15756 12303
rect 15722 12269 15756 12291
rect 15722 12223 15756 12231
rect 15722 12197 15756 12223
rect 15722 12155 15756 12159
rect 15722 12125 15756 12155
rect 15722 12053 15756 12087
rect 15722 11985 15756 12015
rect 15722 11981 15756 11985
rect 15722 11917 15756 11943
rect 15722 11909 15756 11917
rect 15722 11849 15756 11871
rect 15722 11837 15756 11849
rect 15722 11781 15756 11799
rect 15722 11765 15756 11781
rect 15722 11713 15756 11727
rect 15722 11693 15756 11713
rect 15722 11645 15756 11655
rect 15722 11621 15756 11645
rect 15722 11577 15756 11583
rect 15722 11549 15756 11577
rect 15722 11509 15756 11511
rect 15722 11477 15756 11509
rect 15722 11407 15756 11439
rect 15722 11405 15756 11407
rect 15722 11339 15756 11367
rect 15722 11333 15756 11339
rect 15722 11271 15756 11295
rect 15722 11261 15756 11271
rect 15722 11203 15756 11223
rect 15722 11189 15756 11203
rect 15722 11135 15756 11151
rect 15722 11117 15756 11135
rect 15810 13005 15844 13023
rect 15810 12989 15844 13005
rect 15810 12937 15844 12951
rect 15810 12917 15844 12937
rect 15810 12869 15844 12879
rect 15810 12845 15844 12869
rect 15810 12801 15844 12807
rect 15810 12773 15844 12801
rect 15810 12733 15844 12735
rect 15810 12701 15844 12733
rect 15810 12631 15844 12663
rect 15810 12629 15844 12631
rect 15810 12563 15844 12591
rect 15810 12557 15844 12563
rect 15810 12495 15844 12519
rect 15810 12485 15844 12495
rect 15810 12427 15844 12447
rect 15810 12413 15844 12427
rect 15810 12359 15844 12375
rect 15810 12341 15844 12359
rect 15810 12291 15844 12303
rect 15810 12269 15844 12291
rect 15810 12223 15844 12231
rect 15810 12197 15844 12223
rect 15810 12155 15844 12159
rect 15810 12125 15844 12155
rect 15810 12053 15844 12087
rect 15810 11985 15844 12015
rect 15810 11981 15844 11985
rect 15810 11917 15844 11943
rect 15810 11909 15844 11917
rect 15810 11849 15844 11871
rect 15810 11837 15844 11849
rect 15810 11781 15844 11799
rect 15810 11765 15844 11781
rect 15810 11713 15844 11727
rect 15810 11693 15844 11713
rect 15810 11645 15844 11655
rect 15810 11621 15844 11645
rect 15810 11577 15844 11583
rect 15810 11549 15844 11577
rect 15810 11509 15844 11511
rect 15810 11477 15844 11509
rect 15810 11407 15844 11439
rect 15810 11405 15844 11407
rect 15810 11339 15844 11367
rect 15810 11333 15844 11339
rect 15810 11271 15844 11295
rect 15810 11261 15844 11271
rect 15810 11203 15844 11223
rect 15810 11189 15844 11203
rect 15810 11135 15844 11151
rect 15810 11117 15844 11135
rect 15898 13005 15932 13023
rect 15898 12989 15932 13005
rect 15898 12937 15932 12951
rect 15898 12917 15932 12937
rect 15898 12869 15932 12879
rect 15898 12845 15932 12869
rect 15898 12801 15932 12807
rect 15898 12773 15932 12801
rect 15898 12733 15932 12735
rect 15898 12701 15932 12733
rect 15898 12631 15932 12663
rect 15898 12629 15932 12631
rect 15898 12563 15932 12591
rect 15898 12557 15932 12563
rect 15898 12495 15932 12519
rect 15898 12485 15932 12495
rect 15898 12427 15932 12447
rect 15898 12413 15932 12427
rect 15898 12359 15932 12375
rect 15898 12341 15932 12359
rect 15898 12291 15932 12303
rect 15898 12269 15932 12291
rect 15898 12223 15932 12231
rect 15898 12197 15932 12223
rect 15898 12155 15932 12159
rect 15898 12125 15932 12155
rect 15898 12053 15932 12087
rect 15898 11985 15932 12015
rect 15898 11981 15932 11985
rect 15898 11917 15932 11943
rect 15898 11909 15932 11917
rect 15898 11849 15932 11871
rect 15898 11837 15932 11849
rect 15898 11781 15932 11799
rect 15898 11765 15932 11781
rect 15898 11713 15932 11727
rect 15898 11693 15932 11713
rect 15898 11645 15932 11655
rect 15898 11621 15932 11645
rect 15898 11577 15932 11583
rect 15898 11549 15932 11577
rect 15898 11509 15932 11511
rect 15898 11477 15932 11509
rect 15898 11407 15932 11439
rect 15898 11405 15932 11407
rect 15898 11339 15932 11367
rect 15898 11333 15932 11339
rect 15898 11271 15932 11295
rect 15898 11261 15932 11271
rect 15898 11203 15932 11223
rect 15898 11189 15932 11203
rect 15898 11135 15932 11151
rect 15898 11117 15932 11135
rect 15986 13005 16020 13023
rect 15986 12989 16020 13005
rect 15986 12937 16020 12951
rect 15986 12917 16020 12937
rect 15986 12869 16020 12879
rect 15986 12845 16020 12869
rect 15986 12801 16020 12807
rect 15986 12773 16020 12801
rect 15986 12733 16020 12735
rect 15986 12701 16020 12733
rect 15986 12631 16020 12663
rect 15986 12629 16020 12631
rect 15986 12563 16020 12591
rect 15986 12557 16020 12563
rect 15986 12495 16020 12519
rect 15986 12485 16020 12495
rect 15986 12427 16020 12447
rect 15986 12413 16020 12427
rect 15986 12359 16020 12375
rect 15986 12341 16020 12359
rect 15986 12291 16020 12303
rect 15986 12269 16020 12291
rect 15986 12223 16020 12231
rect 15986 12197 16020 12223
rect 15986 12155 16020 12159
rect 15986 12125 16020 12155
rect 15986 12053 16020 12087
rect 15986 11985 16020 12015
rect 15986 11981 16020 11985
rect 15986 11917 16020 11943
rect 15986 11909 16020 11917
rect 15986 11849 16020 11871
rect 15986 11837 16020 11849
rect 15986 11781 16020 11799
rect 15986 11765 16020 11781
rect 15986 11713 16020 11727
rect 15986 11693 16020 11713
rect 15986 11645 16020 11655
rect 15986 11621 16020 11645
rect 15986 11577 16020 11583
rect 15986 11549 16020 11577
rect 15986 11509 16020 11511
rect 15986 11477 16020 11509
rect 15986 11407 16020 11439
rect 15986 11405 16020 11407
rect 15986 11339 16020 11367
rect 15986 11333 16020 11339
rect 15986 11271 16020 11295
rect 15986 11261 16020 11271
rect 15986 11203 16020 11223
rect 15986 11189 16020 11203
rect 15986 11135 16020 11151
rect 15986 11117 16020 11135
rect 16074 13005 16108 13023
rect 16074 12989 16108 13005
rect 16074 12937 16108 12951
rect 16074 12917 16108 12937
rect 16074 12869 16108 12879
rect 16074 12845 16108 12869
rect 16074 12801 16108 12807
rect 16074 12773 16108 12801
rect 16074 12733 16108 12735
rect 16074 12701 16108 12733
rect 16074 12631 16108 12663
rect 16074 12629 16108 12631
rect 16074 12563 16108 12591
rect 16074 12557 16108 12563
rect 16074 12495 16108 12519
rect 16074 12485 16108 12495
rect 16074 12427 16108 12447
rect 16074 12413 16108 12427
rect 16074 12359 16108 12375
rect 16074 12341 16108 12359
rect 16074 12291 16108 12303
rect 16074 12269 16108 12291
rect 16074 12223 16108 12231
rect 16074 12197 16108 12223
rect 16074 12155 16108 12159
rect 16074 12125 16108 12155
rect 16074 12053 16108 12087
rect 16074 11985 16108 12015
rect 16074 11981 16108 11985
rect 16074 11917 16108 11943
rect 16074 11909 16108 11917
rect 16074 11849 16108 11871
rect 16074 11837 16108 11849
rect 16074 11781 16108 11799
rect 16074 11765 16108 11781
rect 16074 11713 16108 11727
rect 16074 11693 16108 11713
rect 16074 11645 16108 11655
rect 16074 11621 16108 11645
rect 16074 11577 16108 11583
rect 16074 11549 16108 11577
rect 16074 11509 16108 11511
rect 16074 11477 16108 11509
rect 16074 11407 16108 11439
rect 16074 11405 16108 11407
rect 16074 11339 16108 11367
rect 16074 11333 16108 11339
rect 16074 11271 16108 11295
rect 16074 11261 16108 11271
rect 16074 11203 16108 11223
rect 16074 11189 16108 11203
rect 16074 11135 16108 11151
rect 16074 11117 16108 11135
rect 16162 13005 16196 13023
rect 16162 12989 16196 13005
rect 16162 12937 16196 12951
rect 16162 12917 16196 12937
rect 16162 12869 16196 12879
rect 16162 12845 16196 12869
rect 16162 12801 16196 12807
rect 16162 12773 16196 12801
rect 16162 12733 16196 12735
rect 16162 12701 16196 12733
rect 16162 12631 16196 12663
rect 16162 12629 16196 12631
rect 16162 12563 16196 12591
rect 16162 12557 16196 12563
rect 16162 12495 16196 12519
rect 16162 12485 16196 12495
rect 16162 12427 16196 12447
rect 16162 12413 16196 12427
rect 16162 12359 16196 12375
rect 16162 12341 16196 12359
rect 16162 12291 16196 12303
rect 16162 12269 16196 12291
rect 16162 12223 16196 12231
rect 16162 12197 16196 12223
rect 16162 12155 16196 12159
rect 16162 12125 16196 12155
rect 16162 12053 16196 12087
rect 16162 11985 16196 12015
rect 16162 11981 16196 11985
rect 16162 11917 16196 11943
rect 16162 11909 16196 11917
rect 16162 11849 16196 11871
rect 16162 11837 16196 11849
rect 16162 11781 16196 11799
rect 16162 11765 16196 11781
rect 16162 11713 16196 11727
rect 16162 11693 16196 11713
rect 16162 11645 16196 11655
rect 16162 11621 16196 11645
rect 16162 11577 16196 11583
rect 16162 11549 16196 11577
rect 16162 11509 16196 11511
rect 16162 11477 16196 11509
rect 16162 11407 16196 11439
rect 16162 11405 16196 11407
rect 16162 11339 16196 11367
rect 16162 11333 16196 11339
rect 16162 11271 16196 11295
rect 16162 11261 16196 11271
rect 16162 11203 16196 11223
rect 16162 11189 16196 11203
rect 16162 11135 16196 11151
rect 16162 11117 16196 11135
rect 16250 13005 16284 13023
rect 16250 12989 16284 13005
rect 16250 12937 16284 12951
rect 16250 12917 16284 12937
rect 16250 12869 16284 12879
rect 16250 12845 16284 12869
rect 16250 12801 16284 12807
rect 16250 12773 16284 12801
rect 16250 12733 16284 12735
rect 16250 12701 16284 12733
rect 16250 12631 16284 12663
rect 16250 12629 16284 12631
rect 16250 12563 16284 12591
rect 16250 12557 16284 12563
rect 16250 12495 16284 12519
rect 16250 12485 16284 12495
rect 16250 12427 16284 12447
rect 16250 12413 16284 12427
rect 16250 12359 16284 12375
rect 16250 12341 16284 12359
rect 16250 12291 16284 12303
rect 16250 12269 16284 12291
rect 16250 12223 16284 12231
rect 16250 12197 16284 12223
rect 16250 12155 16284 12159
rect 16250 12125 16284 12155
rect 16250 12053 16284 12087
rect 16250 11985 16284 12015
rect 16250 11981 16284 11985
rect 16250 11917 16284 11943
rect 16250 11909 16284 11917
rect 16250 11849 16284 11871
rect 16250 11837 16284 11849
rect 16250 11781 16284 11799
rect 16250 11765 16284 11781
rect 16250 11713 16284 11727
rect 16250 11693 16284 11713
rect 16250 11645 16284 11655
rect 16250 11621 16284 11645
rect 16250 11577 16284 11583
rect 16250 11549 16284 11577
rect 16250 11509 16284 11511
rect 16250 11477 16284 11509
rect 16250 11407 16284 11439
rect 16250 11405 16284 11407
rect 16250 11339 16284 11367
rect 16250 11333 16284 11339
rect 16250 11271 16284 11295
rect 16250 11261 16284 11271
rect 16250 11203 16284 11223
rect 16250 11189 16284 11203
rect 16250 11135 16284 11151
rect 16250 11117 16284 11135
rect 16338 13005 16372 13023
rect 16338 12989 16372 13005
rect 16338 12937 16372 12951
rect 16338 12917 16372 12937
rect 16338 12869 16372 12879
rect 16338 12845 16372 12869
rect 16338 12801 16372 12807
rect 16338 12773 16372 12801
rect 16338 12733 16372 12735
rect 16338 12701 16372 12733
rect 16338 12631 16372 12663
rect 16338 12629 16372 12631
rect 16338 12563 16372 12591
rect 16338 12557 16372 12563
rect 16338 12495 16372 12519
rect 16338 12485 16372 12495
rect 16338 12427 16372 12447
rect 16338 12413 16372 12427
rect 16338 12359 16372 12375
rect 16338 12341 16372 12359
rect 16338 12291 16372 12303
rect 16338 12269 16372 12291
rect 16338 12223 16372 12231
rect 16338 12197 16372 12223
rect 16338 12155 16372 12159
rect 16338 12125 16372 12155
rect 16338 12053 16372 12087
rect 16338 11985 16372 12015
rect 16338 11981 16372 11985
rect 16338 11917 16372 11943
rect 16338 11909 16372 11917
rect 16338 11849 16372 11871
rect 16338 11837 16372 11849
rect 16338 11781 16372 11799
rect 16338 11765 16372 11781
rect 16338 11713 16372 11727
rect 16338 11693 16372 11713
rect 16338 11645 16372 11655
rect 16338 11621 16372 11645
rect 16338 11577 16372 11583
rect 16338 11549 16372 11577
rect 16338 11509 16372 11511
rect 16338 11477 16372 11509
rect 16338 11407 16372 11439
rect 16338 11405 16372 11407
rect 16338 11339 16372 11367
rect 16338 11333 16372 11339
rect 16338 11271 16372 11295
rect 16338 11261 16372 11271
rect 16338 11203 16372 11223
rect 16338 11189 16372 11203
rect 16338 11135 16372 11151
rect 16338 11117 16372 11135
rect 16426 13005 16460 13023
rect 16426 12989 16460 13005
rect 16426 12937 16460 12951
rect 16426 12917 16460 12937
rect 16426 12869 16460 12879
rect 16426 12845 16460 12869
rect 16426 12801 16460 12807
rect 16426 12773 16460 12801
rect 16426 12733 16460 12735
rect 16426 12701 16460 12733
rect 16426 12631 16460 12663
rect 16426 12629 16460 12631
rect 16426 12563 16460 12591
rect 16426 12557 16460 12563
rect 16426 12495 16460 12519
rect 16426 12485 16460 12495
rect 16426 12427 16460 12447
rect 16426 12413 16460 12427
rect 16426 12359 16460 12375
rect 16426 12341 16460 12359
rect 16426 12291 16460 12303
rect 16426 12269 16460 12291
rect 16426 12223 16460 12231
rect 16426 12197 16460 12223
rect 16426 12155 16460 12159
rect 16426 12125 16460 12155
rect 16426 12053 16460 12087
rect 16426 11985 16460 12015
rect 16426 11981 16460 11985
rect 16426 11917 16460 11943
rect 16426 11909 16460 11917
rect 16426 11849 16460 11871
rect 16426 11837 16460 11849
rect 16426 11781 16460 11799
rect 16426 11765 16460 11781
rect 16426 11713 16460 11727
rect 16426 11693 16460 11713
rect 16426 11645 16460 11655
rect 16426 11621 16460 11645
rect 16426 11577 16460 11583
rect 16426 11549 16460 11577
rect 16426 11509 16460 11511
rect 16426 11477 16460 11509
rect 16426 11407 16460 11439
rect 16426 11405 16460 11407
rect 16426 11339 16460 11367
rect 16426 11333 16460 11339
rect 16426 11271 16460 11295
rect 16426 11261 16460 11271
rect 16426 11203 16460 11223
rect 16426 11189 16460 11203
rect 16426 11135 16460 11151
rect 16426 11117 16460 11135
rect 16514 13005 16548 13023
rect 16514 12989 16548 13005
rect 16514 12937 16548 12951
rect 16514 12917 16548 12937
rect 16514 12869 16548 12879
rect 16514 12845 16548 12869
rect 16514 12801 16548 12807
rect 16514 12773 16548 12801
rect 16514 12733 16548 12735
rect 16514 12701 16548 12733
rect 16514 12631 16548 12663
rect 16514 12629 16548 12631
rect 16514 12563 16548 12591
rect 16514 12557 16548 12563
rect 16514 12495 16548 12519
rect 16514 12485 16548 12495
rect 16514 12427 16548 12447
rect 16514 12413 16548 12427
rect 16514 12359 16548 12375
rect 16514 12341 16548 12359
rect 16514 12291 16548 12303
rect 16514 12269 16548 12291
rect 16514 12223 16548 12231
rect 16514 12197 16548 12223
rect 16514 12155 16548 12159
rect 16514 12125 16548 12155
rect 16514 12053 16548 12087
rect 16514 11985 16548 12015
rect 16514 11981 16548 11985
rect 16514 11917 16548 11943
rect 16514 11909 16548 11917
rect 16514 11849 16548 11871
rect 16514 11837 16548 11849
rect 16514 11781 16548 11799
rect 16514 11765 16548 11781
rect 16514 11713 16548 11727
rect 16514 11693 16548 11713
rect 16514 11645 16548 11655
rect 16514 11621 16548 11645
rect 16514 11577 16548 11583
rect 16514 11549 16548 11577
rect 16514 11509 16548 11511
rect 16514 11477 16548 11509
rect 16514 11407 16548 11439
rect 16514 11405 16548 11407
rect 16514 11339 16548 11367
rect 16514 11333 16548 11339
rect 16514 11271 16548 11295
rect 16514 11261 16548 11271
rect 16514 11203 16548 11223
rect 16514 11189 16548 11203
rect 16514 11135 16548 11151
rect 16514 11117 16548 11135
rect 16602 13005 16636 13023
rect 16602 12989 16636 13005
rect 16602 12937 16636 12951
rect 16602 12917 16636 12937
rect 16602 12869 16636 12879
rect 16602 12845 16636 12869
rect 16602 12801 16636 12807
rect 16602 12773 16636 12801
rect 16602 12733 16636 12735
rect 16602 12701 16636 12733
rect 16602 12631 16636 12663
rect 16602 12629 16636 12631
rect 16602 12563 16636 12591
rect 16602 12557 16636 12563
rect 16602 12495 16636 12519
rect 16602 12485 16636 12495
rect 16602 12427 16636 12447
rect 16602 12413 16636 12427
rect 16602 12359 16636 12375
rect 16602 12341 16636 12359
rect 16602 12291 16636 12303
rect 16602 12269 16636 12291
rect 16602 12223 16636 12231
rect 16602 12197 16636 12223
rect 16602 12155 16636 12159
rect 16602 12125 16636 12155
rect 16602 12053 16636 12087
rect 16602 11985 16636 12015
rect 16602 11981 16636 11985
rect 16602 11917 16636 11943
rect 16602 11909 16636 11917
rect 16602 11849 16636 11871
rect 16602 11837 16636 11849
rect 16602 11781 16636 11799
rect 16602 11765 16636 11781
rect 16602 11713 16636 11727
rect 16602 11693 16636 11713
rect 16602 11645 16636 11655
rect 16602 11621 16636 11645
rect 16602 11577 16636 11583
rect 16602 11549 16636 11577
rect 16602 11509 16636 11511
rect 16602 11477 16636 11509
rect 16602 11407 16636 11439
rect 16602 11405 16636 11407
rect 16602 11339 16636 11367
rect 16602 11333 16636 11339
rect 16602 11271 16636 11295
rect 16602 11261 16636 11271
rect 16602 11203 16636 11223
rect 16602 11189 16636 11203
rect 16602 11135 16636 11151
rect 16602 11117 16636 11135
rect 16690 13005 16724 13023
rect 16690 12989 16724 13005
rect 16690 12937 16724 12951
rect 16690 12917 16724 12937
rect 16690 12869 16724 12879
rect 16690 12845 16724 12869
rect 16690 12801 16724 12807
rect 16690 12773 16724 12801
rect 16690 12733 16724 12735
rect 16690 12701 16724 12733
rect 16690 12631 16724 12663
rect 16690 12629 16724 12631
rect 16690 12563 16724 12591
rect 16690 12557 16724 12563
rect 16690 12495 16724 12519
rect 16690 12485 16724 12495
rect 16690 12427 16724 12447
rect 16690 12413 16724 12427
rect 16690 12359 16724 12375
rect 16690 12341 16724 12359
rect 16690 12291 16724 12303
rect 16690 12269 16724 12291
rect 16690 12223 16724 12231
rect 16690 12197 16724 12223
rect 16690 12155 16724 12159
rect 16690 12125 16724 12155
rect 16690 12053 16724 12087
rect 16690 11985 16724 12015
rect 16690 11981 16724 11985
rect 16690 11917 16724 11943
rect 16690 11909 16724 11917
rect 16690 11849 16724 11871
rect 16690 11837 16724 11849
rect 16690 11781 16724 11799
rect 16690 11765 16724 11781
rect 16690 11713 16724 11727
rect 16690 11693 16724 11713
rect 16690 11645 16724 11655
rect 16690 11621 16724 11645
rect 16690 11577 16724 11583
rect 16690 11549 16724 11577
rect 16690 11509 16724 11511
rect 16690 11477 16724 11509
rect 16690 11407 16724 11439
rect 16690 11405 16724 11407
rect 16690 11339 16724 11367
rect 16690 11333 16724 11339
rect 16690 11271 16724 11295
rect 16690 11261 16724 11271
rect 16690 11203 16724 11223
rect 16690 11189 16724 11203
rect 16690 11135 16724 11151
rect 16690 11117 16724 11135
rect 16778 13005 16812 13023
rect 16778 12989 16812 13005
rect 16778 12937 16812 12951
rect 16778 12917 16812 12937
rect 16778 12869 16812 12879
rect 16778 12845 16812 12869
rect 16778 12801 16812 12807
rect 16778 12773 16812 12801
rect 16778 12733 16812 12735
rect 16778 12701 16812 12733
rect 16778 12631 16812 12663
rect 16778 12629 16812 12631
rect 16778 12563 16812 12591
rect 16778 12557 16812 12563
rect 16778 12495 16812 12519
rect 16778 12485 16812 12495
rect 16778 12427 16812 12447
rect 16778 12413 16812 12427
rect 16778 12359 16812 12375
rect 16778 12341 16812 12359
rect 16778 12291 16812 12303
rect 16778 12269 16812 12291
rect 16778 12223 16812 12231
rect 16778 12197 16812 12223
rect 16778 12155 16812 12159
rect 16778 12125 16812 12155
rect 16778 12053 16812 12087
rect 16778 11985 16812 12015
rect 16778 11981 16812 11985
rect 16778 11917 16812 11943
rect 16778 11909 16812 11917
rect 16778 11849 16812 11871
rect 16778 11837 16812 11849
rect 16778 11781 16812 11799
rect 16778 11765 16812 11781
rect 16778 11713 16812 11727
rect 16778 11693 16812 11713
rect 16778 11645 16812 11655
rect 16778 11621 16812 11645
rect 16778 11577 16812 11583
rect 16778 11549 16812 11577
rect 16778 11509 16812 11511
rect 16778 11477 16812 11509
rect 16778 11407 16812 11439
rect 16778 11405 16812 11407
rect 16778 11339 16812 11367
rect 16778 11333 16812 11339
rect 16778 11271 16812 11295
rect 16778 11261 16812 11271
rect 16778 11203 16812 11223
rect 16778 11189 16812 11203
rect 16778 11135 16812 11151
rect 16778 11117 16812 11135
rect 16866 13005 16900 13023
rect 16866 12989 16900 13005
rect 16866 12937 16900 12951
rect 16866 12917 16900 12937
rect 16866 12869 16900 12879
rect 16866 12845 16900 12869
rect 16866 12801 16900 12807
rect 16866 12773 16900 12801
rect 16866 12733 16900 12735
rect 16866 12701 16900 12733
rect 16866 12631 16900 12663
rect 16866 12629 16900 12631
rect 16866 12563 16900 12591
rect 16866 12557 16900 12563
rect 16866 12495 16900 12519
rect 16866 12485 16900 12495
rect 16866 12427 16900 12447
rect 16866 12413 16900 12427
rect 16866 12359 16900 12375
rect 16866 12341 16900 12359
rect 16866 12291 16900 12303
rect 16866 12269 16900 12291
rect 16866 12223 16900 12231
rect 16866 12197 16900 12223
rect 16866 12155 16900 12159
rect 16866 12125 16900 12155
rect 16866 12053 16900 12087
rect 16866 11985 16900 12015
rect 16866 11981 16900 11985
rect 16866 11917 16900 11943
rect 16866 11909 16900 11917
rect 16866 11849 16900 11871
rect 16866 11837 16900 11849
rect 16866 11781 16900 11799
rect 16866 11765 16900 11781
rect 16866 11713 16900 11727
rect 16866 11693 16900 11713
rect 16866 11645 16900 11655
rect 16866 11621 16900 11645
rect 16866 11577 16900 11583
rect 16866 11549 16900 11577
rect 16866 11509 16900 11511
rect 16866 11477 16900 11509
rect 16866 11407 16900 11439
rect 16866 11405 16900 11407
rect 16866 11339 16900 11367
rect 16866 11333 16900 11339
rect 16866 11271 16900 11295
rect 16866 11261 16900 11271
rect 16866 11203 16900 11223
rect 16866 11189 16900 11203
rect 16866 11135 16900 11151
rect 16866 11117 16900 11135
rect 16954 13005 16988 13023
rect 16954 12989 16988 13005
rect 16954 12937 16988 12951
rect 16954 12917 16988 12937
rect 16954 12869 16988 12879
rect 16954 12845 16988 12869
rect 16954 12801 16988 12807
rect 16954 12773 16988 12801
rect 16954 12733 16988 12735
rect 16954 12701 16988 12733
rect 16954 12631 16988 12663
rect 16954 12629 16988 12631
rect 16954 12563 16988 12591
rect 16954 12557 16988 12563
rect 16954 12495 16988 12519
rect 16954 12485 16988 12495
rect 16954 12427 16988 12447
rect 16954 12413 16988 12427
rect 16954 12359 16988 12375
rect 16954 12341 16988 12359
rect 16954 12291 16988 12303
rect 16954 12269 16988 12291
rect 16954 12223 16988 12231
rect 16954 12197 16988 12223
rect 16954 12155 16988 12159
rect 16954 12125 16988 12155
rect 16954 12053 16988 12087
rect 16954 11985 16988 12015
rect 16954 11981 16988 11985
rect 16954 11917 16988 11943
rect 16954 11909 16988 11917
rect 16954 11849 16988 11871
rect 16954 11837 16988 11849
rect 16954 11781 16988 11799
rect 16954 11765 16988 11781
rect 16954 11713 16988 11727
rect 16954 11693 16988 11713
rect 16954 11645 16988 11655
rect 16954 11621 16988 11645
rect 16954 11577 16988 11583
rect 16954 11549 16988 11577
rect 16954 11509 16988 11511
rect 16954 11477 16988 11509
rect 16954 11407 16988 11439
rect 16954 11405 16988 11407
rect 16954 11339 16988 11367
rect 16954 11333 16988 11339
rect 16954 11271 16988 11295
rect 16954 11261 16988 11271
rect 16954 11203 16988 11223
rect 16954 11189 16988 11203
rect 16954 11135 16988 11151
rect 16954 11117 16988 11135
rect 17042 13005 17076 13023
rect 17042 12989 17076 13005
rect 17042 12937 17076 12951
rect 17042 12917 17076 12937
rect 17042 12869 17076 12879
rect 17042 12845 17076 12869
rect 17042 12801 17076 12807
rect 17042 12773 17076 12801
rect 17042 12733 17076 12735
rect 17042 12701 17076 12733
rect 17042 12631 17076 12663
rect 17042 12629 17076 12631
rect 17042 12563 17076 12591
rect 17042 12557 17076 12563
rect 17042 12495 17076 12519
rect 17042 12485 17076 12495
rect 17042 12427 17076 12447
rect 17042 12413 17076 12427
rect 17042 12359 17076 12375
rect 17042 12341 17076 12359
rect 17042 12291 17076 12303
rect 17042 12269 17076 12291
rect 17042 12223 17076 12231
rect 17042 12197 17076 12223
rect 17042 12155 17076 12159
rect 17042 12125 17076 12155
rect 17042 12053 17076 12087
rect 17042 11985 17076 12015
rect 17042 11981 17076 11985
rect 17042 11917 17076 11943
rect 17042 11909 17076 11917
rect 17042 11849 17076 11871
rect 17042 11837 17076 11849
rect 17042 11781 17076 11799
rect 17042 11765 17076 11781
rect 17042 11713 17076 11727
rect 17042 11693 17076 11713
rect 17042 11645 17076 11655
rect 17042 11621 17076 11645
rect 17042 11577 17076 11583
rect 17042 11549 17076 11577
rect 17042 11509 17076 11511
rect 17042 11477 17076 11509
rect 17042 11407 17076 11439
rect 17042 11405 17076 11407
rect 17042 11339 17076 11367
rect 17042 11333 17076 11339
rect 17042 11271 17076 11295
rect 17042 11261 17076 11271
rect 17042 11203 17076 11223
rect 17042 11189 17076 11203
rect 17042 11135 17076 11151
rect 17042 11117 17076 11135
rect 17130 13005 17164 13023
rect 17130 12989 17164 13005
rect 17130 12937 17164 12951
rect 17130 12917 17164 12937
rect 17130 12869 17164 12879
rect 17130 12845 17164 12869
rect 17130 12801 17164 12807
rect 17130 12773 17164 12801
rect 17130 12733 17164 12735
rect 17130 12701 17164 12733
rect 17130 12631 17164 12663
rect 17130 12629 17164 12631
rect 17130 12563 17164 12591
rect 17130 12557 17164 12563
rect 17130 12495 17164 12519
rect 17130 12485 17164 12495
rect 17130 12427 17164 12447
rect 17130 12413 17164 12427
rect 17130 12359 17164 12375
rect 17130 12341 17164 12359
rect 17130 12291 17164 12303
rect 17130 12269 17164 12291
rect 17130 12223 17164 12231
rect 17130 12197 17164 12223
rect 17130 12155 17164 12159
rect 17130 12125 17164 12155
rect 17130 12053 17164 12087
rect 17130 11985 17164 12015
rect 17130 11981 17164 11985
rect 17130 11917 17164 11943
rect 17130 11909 17164 11917
rect 17130 11849 17164 11871
rect 17130 11837 17164 11849
rect 17130 11781 17164 11799
rect 17130 11765 17164 11781
rect 17130 11713 17164 11727
rect 17130 11693 17164 11713
rect 17130 11645 17164 11655
rect 17130 11621 17164 11645
rect 17130 11577 17164 11583
rect 17130 11549 17164 11577
rect 17130 11509 17164 11511
rect 17130 11477 17164 11509
rect 17130 11407 17164 11439
rect 17130 11405 17164 11407
rect 17130 11339 17164 11367
rect 17130 11333 17164 11339
rect 17130 11271 17164 11295
rect 17130 11261 17164 11271
rect 17130 11203 17164 11223
rect 17130 11189 17164 11203
rect 17130 11135 17164 11151
rect 17130 11117 17164 11135
rect 17218 13005 17252 13023
rect 17218 12989 17252 13005
rect 17218 12937 17252 12951
rect 17218 12917 17252 12937
rect 17218 12869 17252 12879
rect 17218 12845 17252 12869
rect 17218 12801 17252 12807
rect 17218 12773 17252 12801
rect 17218 12733 17252 12735
rect 17218 12701 17252 12733
rect 17218 12631 17252 12663
rect 17218 12629 17252 12631
rect 17218 12563 17252 12591
rect 17218 12557 17252 12563
rect 17218 12495 17252 12519
rect 17218 12485 17252 12495
rect 17218 12427 17252 12447
rect 17218 12413 17252 12427
rect 17218 12359 17252 12375
rect 17218 12341 17252 12359
rect 17218 12291 17252 12303
rect 17218 12269 17252 12291
rect 17218 12223 17252 12231
rect 17218 12197 17252 12223
rect 17218 12155 17252 12159
rect 17218 12125 17252 12155
rect 17218 12053 17252 12087
rect 17218 11985 17252 12015
rect 17218 11981 17252 11985
rect 17218 11917 17252 11943
rect 17218 11909 17252 11917
rect 17218 11849 17252 11871
rect 17218 11837 17252 11849
rect 17218 11781 17252 11799
rect 17218 11765 17252 11781
rect 17218 11713 17252 11727
rect 17218 11693 17252 11713
rect 17218 11645 17252 11655
rect 17218 11621 17252 11645
rect 17218 11577 17252 11583
rect 17218 11549 17252 11577
rect 17218 11509 17252 11511
rect 17218 11477 17252 11509
rect 17218 11407 17252 11439
rect 17218 11405 17252 11407
rect 17218 11339 17252 11367
rect 17218 11333 17252 11339
rect 17218 11271 17252 11295
rect 17218 11261 17252 11271
rect 17218 11203 17252 11223
rect 17218 11189 17252 11203
rect 17218 11135 17252 11151
rect 17218 11117 17252 11135
rect 17306 13005 17340 13023
rect 17306 12989 17340 13005
rect 17306 12937 17340 12951
rect 17306 12917 17340 12937
rect 17306 12869 17340 12879
rect 17306 12845 17340 12869
rect 17306 12801 17340 12807
rect 17306 12773 17340 12801
rect 17306 12733 17340 12735
rect 17306 12701 17340 12733
rect 17306 12631 17340 12663
rect 17306 12629 17340 12631
rect 17306 12563 17340 12591
rect 17306 12557 17340 12563
rect 17306 12495 17340 12519
rect 17306 12485 17340 12495
rect 17306 12427 17340 12447
rect 17306 12413 17340 12427
rect 17306 12359 17340 12375
rect 17306 12341 17340 12359
rect 17306 12291 17340 12303
rect 17306 12269 17340 12291
rect 17306 12223 17340 12231
rect 17306 12197 17340 12223
rect 17306 12155 17340 12159
rect 17306 12125 17340 12155
rect 17306 12053 17340 12087
rect 17306 11985 17340 12015
rect 17306 11981 17340 11985
rect 17306 11917 17340 11943
rect 17306 11909 17340 11917
rect 17306 11849 17340 11871
rect 17306 11837 17340 11849
rect 17306 11781 17340 11799
rect 17306 11765 17340 11781
rect 17306 11713 17340 11727
rect 17306 11693 17340 11713
rect 17306 11645 17340 11655
rect 17306 11621 17340 11645
rect 17306 11577 17340 11583
rect 17306 11549 17340 11577
rect 17306 11509 17340 11511
rect 17306 11477 17340 11509
rect 17306 11407 17340 11439
rect 17306 11405 17340 11407
rect 17306 11339 17340 11367
rect 17306 11333 17340 11339
rect 17306 11271 17340 11295
rect 17306 11261 17340 11271
rect 17306 11203 17340 11223
rect 17306 11189 17340 11203
rect 17306 11135 17340 11151
rect 17306 11117 17340 11135
rect 17394 13005 17428 13023
rect 17394 12989 17428 13005
rect 17394 12937 17428 12951
rect 17394 12917 17428 12937
rect 17394 12869 17428 12879
rect 17394 12845 17428 12869
rect 17394 12801 17428 12807
rect 17394 12773 17428 12801
rect 17394 12733 17428 12735
rect 17394 12701 17428 12733
rect 17394 12631 17428 12663
rect 17394 12629 17428 12631
rect 17394 12563 17428 12591
rect 17394 12557 17428 12563
rect 17394 12495 17428 12519
rect 17394 12485 17428 12495
rect 17394 12427 17428 12447
rect 17394 12413 17428 12427
rect 17394 12359 17428 12375
rect 17394 12341 17428 12359
rect 17394 12291 17428 12303
rect 17394 12269 17428 12291
rect 17394 12223 17428 12231
rect 17394 12197 17428 12223
rect 17394 12155 17428 12159
rect 17394 12125 17428 12155
rect 17394 12053 17428 12087
rect 17394 11985 17428 12015
rect 17394 11981 17428 11985
rect 17394 11917 17428 11943
rect 17394 11909 17428 11917
rect 17394 11849 17428 11871
rect 17394 11837 17428 11849
rect 17394 11781 17428 11799
rect 17394 11765 17428 11781
rect 17394 11713 17428 11727
rect 17394 11693 17428 11713
rect 17394 11645 17428 11655
rect 17394 11621 17428 11645
rect 17394 11577 17428 11583
rect 17394 11549 17428 11577
rect 17394 11509 17428 11511
rect 17394 11477 17428 11509
rect 17394 11407 17428 11439
rect 17394 11405 17428 11407
rect 17394 11339 17428 11367
rect 17394 11333 17428 11339
rect 17394 11271 17428 11295
rect 17394 11261 17428 11271
rect 17394 11203 17428 11223
rect 17394 11189 17428 11203
rect 17394 11135 17428 11151
rect 17394 11117 17428 11135
rect 17482 13005 17516 13023
rect 17482 12989 17516 13005
rect 17482 12937 17516 12951
rect 17482 12917 17516 12937
rect 17482 12869 17516 12879
rect 17482 12845 17516 12869
rect 17482 12801 17516 12807
rect 17482 12773 17516 12801
rect 17482 12733 17516 12735
rect 17482 12701 17516 12733
rect 17482 12631 17516 12663
rect 17482 12629 17516 12631
rect 17482 12563 17516 12591
rect 17482 12557 17516 12563
rect 17482 12495 17516 12519
rect 17482 12485 17516 12495
rect 17482 12427 17516 12447
rect 17482 12413 17516 12427
rect 17482 12359 17516 12375
rect 17482 12341 17516 12359
rect 17482 12291 17516 12303
rect 17482 12269 17516 12291
rect 17482 12223 17516 12231
rect 17482 12197 17516 12223
rect 17482 12155 17516 12159
rect 17482 12125 17516 12155
rect 17482 12053 17516 12087
rect 17482 11985 17516 12015
rect 17482 11981 17516 11985
rect 17482 11917 17516 11943
rect 17482 11909 17516 11917
rect 17482 11849 17516 11871
rect 17482 11837 17516 11849
rect 17482 11781 17516 11799
rect 17482 11765 17516 11781
rect 17482 11713 17516 11727
rect 17482 11693 17516 11713
rect 17482 11645 17516 11655
rect 17482 11621 17516 11645
rect 17482 11577 17516 11583
rect 17482 11549 17516 11577
rect 17482 11509 17516 11511
rect 17482 11477 17516 11509
rect 17482 11407 17516 11439
rect 17482 11405 17516 11407
rect 17482 11339 17516 11367
rect 17482 11333 17516 11339
rect 17482 11271 17516 11295
rect 17482 11261 17516 11271
rect 17482 11203 17516 11223
rect 17482 11189 17516 11203
rect 17482 11135 17516 11151
rect 17482 11117 17516 11135
rect 13514 10827 13548 10861
rect 17395 10812 17429 10846
rect 14503 10693 14537 10701
rect 14575 10693 14609 10701
rect 14647 10693 14681 10701
rect 14503 10667 14527 10693
rect 14527 10667 14537 10693
rect 14575 10667 14595 10693
rect 14595 10667 14609 10693
rect 14647 10667 14663 10693
rect 14663 10667 14681 10693
rect 13929 8972 16915 9654
<< metal1 >>
rect 2229 28863 28685 28930
rect 2229 28815 27191 28863
rect 2229 28791 14128 28815
rect 2229 27715 2351 28791
rect 3683 27715 14128 28791
rect 2229 27701 14128 27715
rect 16394 27787 27191 28815
rect 28523 27787 28685 28863
rect 16394 27701 28685 27787
rect 2229 27600 28685 27701
rect 4162 26936 26614 26978
rect 4162 26928 25306 26936
rect 4162 25660 4248 26928
rect 5516 25668 25306 26928
rect 26574 25668 26614 26936
rect 5516 25660 26614 25668
rect 4162 25554 26614 25660
rect 16810 24606 16910 24620
rect 13052 24598 13473 24606
rect 13052 24564 13065 24598
rect 13099 24564 13137 24598
rect 13171 24564 13209 24598
rect 13243 24564 13281 24598
rect 13315 24564 13353 24598
rect 13387 24564 13425 24598
rect 13459 24564 13473 24598
rect 13052 24556 13473 24564
rect 16483 24598 16910 24606
rect 16483 24564 16496 24598
rect 16530 24564 16568 24598
rect 16602 24564 16640 24598
rect 16674 24564 16712 24598
rect 16746 24564 16784 24598
rect 16818 24591 16856 24598
rect 16818 24564 16834 24591
rect 16890 24564 16910 24598
rect 16483 24556 16834 24564
rect 16810 24539 16834 24556
rect 16886 24539 16910 24564
rect 16810 24510 16910 24539
rect 12535 24142 16435 24280
rect 12535 24140 16441 24142
rect 12535 24112 17620 24140
rect 12535 24078 16806 24112
rect 16840 24078 16998 24112
rect 17032 24078 17190 24112
rect 17224 24078 17382 24112
rect 17416 24078 17574 24112
rect 17608 24078 17620 24112
rect 12535 24070 17620 24078
rect 12535 24003 16441 24070
rect 12535 17956 12812 24003
rect 13070 23926 13340 23940
rect 13070 23918 13503 23926
rect 13070 23884 13095 23918
rect 13129 23884 13167 23918
rect 13201 23884 13239 23918
rect 13273 23884 13311 23918
rect 13345 23884 13383 23918
rect 13417 23884 13455 23918
rect 13489 23884 13503 23918
rect 13070 23876 13503 23884
rect 14303 23918 16441 24003
rect 14303 23884 14326 23918
rect 14360 23884 14398 23918
rect 14432 23884 14470 23918
rect 14504 23884 14542 23918
rect 14576 23884 14614 23918
rect 14648 23884 14686 23918
rect 14720 23884 16441 23918
rect 13070 23523 13340 23876
rect 14303 23865 16441 23884
rect 16656 23993 16702 24040
rect 16656 23959 16662 23993
rect 16696 23959 16702 23993
rect 16656 23921 16702 23959
rect 16656 23887 16662 23921
rect 16696 23887 16702 23921
rect 16743 24001 16813 24041
rect 16743 23949 16750 24001
rect 16802 23949 16813 24001
rect 16743 23921 16813 23949
rect 16743 23911 16758 23921
rect 16656 23849 16702 23887
rect 16656 23815 16662 23849
rect 16696 23815 16702 23849
rect 16656 23777 16702 23815
rect 16656 23743 16662 23777
rect 16696 23743 16702 23777
rect 16656 23705 16702 23743
rect 16656 23671 16662 23705
rect 16696 23671 16702 23705
rect 16656 23633 16702 23671
rect 13070 23417 13111 23523
rect 13289 23417 13340 23523
rect 13070 23370 13340 23417
rect 15260 23610 15432 23632
rect 13648 23361 13802 23388
rect 13648 23053 13670 23361
rect 13786 23053 13802 23361
rect 15260 23366 15285 23610
rect 15401 23366 15432 23610
rect 16656 23599 16662 23633
rect 16696 23599 16702 23633
rect 16270 23553 16450 23580
rect 16270 23437 16302 23553
rect 16418 23437 16450 23553
rect 16270 23410 16450 23437
rect 16656 23561 16702 23599
rect 16656 23527 16662 23561
rect 16696 23527 16702 23561
rect 16656 23489 16702 23527
rect 16656 23455 16662 23489
rect 16696 23455 16702 23489
rect 16656 23417 16702 23455
rect 15260 23312 15432 23366
rect 16656 23383 16662 23417
rect 16696 23383 16702 23417
rect 16656 23345 16702 23383
rect 14090 23222 14740 23240
rect 14090 23188 14114 23222
rect 14148 23188 14306 23222
rect 14340 23188 14498 23222
rect 14532 23188 14690 23222
rect 14724 23188 14740 23222
rect 14090 23180 14740 23188
rect 15260 23210 15420 23312
rect 16656 23311 16662 23345
rect 16696 23311 16702 23345
rect 15950 23270 16030 23280
rect 15950 23236 15974 23270
rect 16008 23236 16030 23270
rect 15950 23230 16030 23236
rect 16656 23273 16702 23311
rect 16656 23239 16662 23273
rect 16696 23239 16702 23273
rect 15260 23176 15324 23210
rect 15358 23176 15420 23210
rect 16656 23201 16702 23239
rect 13648 23028 13802 23053
rect 13964 23103 14010 23150
rect 13964 23069 13970 23103
rect 14004 23069 14010 23103
rect 13964 23031 14010 23069
rect 14041 23117 14111 23151
rect 14041 23065 14050 23117
rect 14102 23065 14111 23117
rect 14041 23031 14111 23065
rect 14156 23103 14202 23150
rect 14156 23069 14162 23103
rect 14196 23069 14202 23103
rect 14156 23031 14202 23069
rect 14241 23117 14311 23151
rect 14241 23065 14250 23117
rect 14302 23065 14311 23117
rect 14241 23031 14311 23065
rect 14348 23103 14394 23150
rect 14348 23069 14354 23103
rect 14388 23069 14394 23103
rect 14348 23031 14394 23069
rect 14431 23117 14501 23151
rect 14431 23065 14440 23117
rect 14492 23065 14501 23117
rect 14431 23031 14501 23065
rect 14540 23103 14586 23150
rect 14540 23069 14546 23103
rect 14580 23069 14586 23103
rect 14540 23031 14586 23069
rect 14621 23117 14691 23151
rect 14621 23065 14630 23117
rect 14682 23065 14691 23117
rect 14621 23031 14691 23065
rect 14732 23103 14778 23150
rect 14732 23069 14738 23103
rect 14772 23069 14778 23103
rect 14732 23031 14778 23069
rect 13496 22050 13546 22064
rect 13496 22016 13504 22050
rect 13538 22016 13546 22050
rect 13496 21978 13546 22016
rect 13496 21944 13504 21978
rect 13538 21944 13546 21978
rect 13496 21906 13546 21944
rect 13496 21872 13504 21906
rect 13538 21872 13546 21906
rect 13496 21834 13546 21872
rect 13496 21800 13504 21834
rect 13538 21800 13546 21834
rect 13496 21780 13546 21800
rect 13650 21780 13800 23028
rect 13480 21762 13800 21780
rect 13480 21728 13504 21762
rect 13538 21728 13800 21762
rect 13480 21690 13800 21728
rect 13480 21656 13504 21690
rect 13538 21656 13800 21690
rect 13480 21630 13800 21656
rect 13496 21519 13546 21533
rect 13496 21485 13504 21519
rect 13538 21485 13546 21519
rect 13496 21447 13546 21485
rect 13496 21413 13504 21447
rect 13538 21413 13546 21447
rect 13496 21375 13546 21413
rect 13496 21341 13504 21375
rect 13538 21341 13546 21375
rect 13496 21303 13546 21341
rect 13496 21269 13504 21303
rect 13538 21269 13546 21303
rect 13496 21231 13546 21269
rect 13496 21197 13504 21231
rect 13538 21197 13546 21231
rect 13496 21190 13546 21197
rect 12535 17712 12585 17956
rect 12765 17712 12812 17956
rect 12535 17676 12812 17712
rect 13000 21159 13560 21190
rect 13000 21125 13504 21159
rect 13538 21125 13560 21159
rect 13000 21070 13560 21125
rect 13710 21120 13800 21630
rect 13964 22997 13970 23031
rect 14004 22997 14010 23031
rect 13964 22959 14010 22997
rect 13964 22925 13970 22959
rect 14004 22925 14010 22959
rect 13964 22887 14010 22925
rect 13964 22853 13970 22887
rect 14004 22853 14010 22887
rect 13964 22815 14010 22853
rect 13964 22781 13970 22815
rect 14004 22781 14010 22815
rect 13964 22743 14010 22781
rect 13964 22709 13970 22743
rect 14004 22709 14010 22743
rect 13964 22671 14010 22709
rect 13964 22637 13970 22671
rect 14004 22637 14010 22671
rect 13964 22599 14010 22637
rect 13964 22565 13970 22599
rect 14004 22565 14010 22599
rect 13964 22527 14010 22565
rect 13964 22493 13970 22527
rect 14004 22493 14010 22527
rect 13964 22455 14010 22493
rect 13964 22421 13970 22455
rect 14004 22421 14010 22455
rect 13964 22383 14010 22421
rect 13964 22349 13970 22383
rect 14004 22349 14010 22383
rect 13964 22311 14010 22349
rect 13964 22277 13970 22311
rect 14004 22277 14010 22311
rect 13964 22239 14010 22277
rect 13964 22205 13970 22239
rect 14004 22205 14010 22239
rect 13964 22167 14010 22205
rect 13964 22133 13970 22167
rect 14004 22133 14010 22167
rect 13964 22095 14010 22133
rect 13964 22061 13970 22095
rect 14004 22061 14010 22095
rect 13964 22023 14010 22061
rect 13964 21989 13970 22023
rect 14004 21989 14010 22023
rect 13964 21951 14010 21989
rect 13964 21917 13970 21951
rect 14004 21917 14010 21951
rect 13964 21879 14010 21917
rect 13964 21845 13970 21879
rect 14004 21845 14010 21879
rect 13964 21807 14010 21845
rect 13964 21773 13970 21807
rect 14004 21773 14010 21807
rect 13964 21735 14010 21773
rect 13964 21701 13970 21735
rect 14004 21701 14010 21735
rect 13964 21663 14010 21701
rect 13964 21629 13970 21663
rect 14004 21629 14010 21663
rect 13964 21591 14010 21629
rect 13964 21557 13970 21591
rect 14004 21557 14010 21591
rect 13964 21519 14010 21557
rect 13964 21485 13970 21519
rect 14004 21485 14010 21519
rect 13964 21447 14010 21485
rect 13964 21413 13970 21447
rect 14004 21413 14010 21447
rect 13964 21375 14010 21413
rect 13964 21341 13970 21375
rect 14004 21341 14010 21375
rect 13964 21303 14010 21341
rect 13964 21271 13970 21303
rect 13951 21269 13970 21271
rect 14004 21271 14010 21303
rect 14060 22997 14066 23031
rect 14100 22997 14106 23031
rect 14060 22959 14106 22997
rect 14060 22925 14066 22959
rect 14100 22925 14106 22959
rect 14060 22887 14106 22925
rect 14060 22853 14066 22887
rect 14100 22853 14106 22887
rect 14060 22815 14106 22853
rect 14060 22781 14066 22815
rect 14100 22781 14106 22815
rect 14060 22743 14106 22781
rect 14060 22709 14066 22743
rect 14100 22709 14106 22743
rect 14060 22671 14106 22709
rect 14060 22637 14066 22671
rect 14100 22637 14106 22671
rect 14060 22599 14106 22637
rect 14060 22565 14066 22599
rect 14100 22565 14106 22599
rect 14060 22527 14106 22565
rect 14060 22493 14066 22527
rect 14100 22493 14106 22527
rect 14060 22455 14106 22493
rect 14060 22421 14066 22455
rect 14100 22421 14106 22455
rect 14060 22383 14106 22421
rect 14060 22349 14066 22383
rect 14100 22349 14106 22383
rect 14060 22311 14106 22349
rect 14060 22277 14066 22311
rect 14100 22277 14106 22311
rect 14060 22239 14106 22277
rect 14060 22205 14066 22239
rect 14100 22205 14106 22239
rect 14060 22167 14106 22205
rect 14060 22133 14066 22167
rect 14100 22133 14106 22167
rect 14060 22095 14106 22133
rect 14060 22061 14066 22095
rect 14100 22061 14106 22095
rect 14060 22023 14106 22061
rect 14060 21989 14066 22023
rect 14100 21989 14106 22023
rect 14060 21951 14106 21989
rect 14060 21917 14066 21951
rect 14100 21917 14106 21951
rect 14060 21879 14106 21917
rect 14060 21845 14066 21879
rect 14100 21845 14106 21879
rect 14060 21807 14106 21845
rect 14060 21773 14066 21807
rect 14100 21773 14106 21807
rect 14060 21735 14106 21773
rect 14060 21701 14066 21735
rect 14100 21701 14106 21735
rect 14060 21663 14106 21701
rect 14060 21629 14066 21663
rect 14100 21629 14106 21663
rect 14060 21591 14106 21629
rect 14060 21557 14066 21591
rect 14100 21557 14106 21591
rect 14060 21519 14106 21557
rect 14060 21485 14066 21519
rect 14100 21485 14106 21519
rect 14060 21447 14106 21485
rect 14060 21413 14066 21447
rect 14100 21413 14106 21447
rect 14060 21375 14106 21413
rect 14060 21341 14066 21375
rect 14100 21341 14106 21375
rect 14060 21303 14106 21341
rect 14004 21269 14021 21271
rect 13951 21237 14021 21269
rect 13951 21185 13960 21237
rect 14012 21185 14021 21237
rect 13951 21151 14021 21185
rect 14060 21269 14066 21303
rect 14100 21269 14106 21303
rect 14156 22997 14162 23031
rect 14196 22997 14202 23031
rect 14156 22959 14202 22997
rect 14156 22925 14162 22959
rect 14196 22925 14202 22959
rect 14156 22887 14202 22925
rect 14156 22853 14162 22887
rect 14196 22853 14202 22887
rect 14156 22815 14202 22853
rect 14156 22781 14162 22815
rect 14196 22781 14202 22815
rect 14156 22743 14202 22781
rect 14156 22709 14162 22743
rect 14196 22709 14202 22743
rect 14156 22671 14202 22709
rect 14156 22637 14162 22671
rect 14196 22637 14202 22671
rect 14156 22599 14202 22637
rect 14156 22565 14162 22599
rect 14196 22565 14202 22599
rect 14156 22527 14202 22565
rect 14156 22493 14162 22527
rect 14196 22493 14202 22527
rect 14156 22455 14202 22493
rect 14156 22421 14162 22455
rect 14196 22421 14202 22455
rect 14156 22383 14202 22421
rect 14156 22349 14162 22383
rect 14196 22349 14202 22383
rect 14156 22311 14202 22349
rect 14156 22277 14162 22311
rect 14196 22277 14202 22311
rect 14156 22239 14202 22277
rect 14156 22205 14162 22239
rect 14196 22205 14202 22239
rect 14156 22167 14202 22205
rect 14156 22133 14162 22167
rect 14196 22133 14202 22167
rect 14156 22095 14202 22133
rect 14156 22061 14162 22095
rect 14196 22061 14202 22095
rect 14156 22023 14202 22061
rect 14156 21989 14162 22023
rect 14196 21989 14202 22023
rect 14156 21951 14202 21989
rect 14156 21917 14162 21951
rect 14196 21917 14202 21951
rect 14156 21879 14202 21917
rect 14156 21845 14162 21879
rect 14196 21845 14202 21879
rect 14156 21807 14202 21845
rect 14156 21773 14162 21807
rect 14196 21773 14202 21807
rect 14156 21735 14202 21773
rect 14156 21701 14162 21735
rect 14196 21701 14202 21735
rect 14156 21663 14202 21701
rect 14156 21629 14162 21663
rect 14196 21629 14202 21663
rect 14156 21591 14202 21629
rect 14156 21557 14162 21591
rect 14196 21557 14202 21591
rect 14156 21519 14202 21557
rect 14156 21485 14162 21519
rect 14196 21485 14202 21519
rect 14156 21447 14202 21485
rect 14156 21413 14162 21447
rect 14196 21413 14202 21447
rect 14156 21375 14202 21413
rect 14156 21341 14162 21375
rect 14196 21341 14202 21375
rect 14156 21303 14202 21341
rect 14156 21271 14162 21303
rect 14060 21231 14106 21269
rect 14060 21197 14066 21231
rect 14100 21197 14106 21231
rect 13964 21150 14010 21151
rect 14060 21150 14106 21197
rect 14141 21269 14162 21271
rect 14196 21271 14202 21303
rect 14252 22997 14258 23031
rect 14292 22997 14298 23031
rect 14252 22959 14298 22997
rect 14252 22925 14258 22959
rect 14292 22925 14298 22959
rect 14252 22887 14298 22925
rect 14252 22853 14258 22887
rect 14292 22853 14298 22887
rect 14252 22815 14298 22853
rect 14252 22781 14258 22815
rect 14292 22781 14298 22815
rect 14252 22743 14298 22781
rect 14252 22709 14258 22743
rect 14292 22709 14298 22743
rect 14252 22671 14298 22709
rect 14252 22637 14258 22671
rect 14292 22637 14298 22671
rect 14252 22599 14298 22637
rect 14252 22565 14258 22599
rect 14292 22565 14298 22599
rect 14252 22527 14298 22565
rect 14252 22493 14258 22527
rect 14292 22493 14298 22527
rect 14252 22455 14298 22493
rect 14252 22421 14258 22455
rect 14292 22421 14298 22455
rect 14252 22383 14298 22421
rect 14252 22349 14258 22383
rect 14292 22349 14298 22383
rect 14252 22311 14298 22349
rect 14252 22277 14258 22311
rect 14292 22277 14298 22311
rect 14252 22239 14298 22277
rect 14252 22205 14258 22239
rect 14292 22205 14298 22239
rect 14252 22167 14298 22205
rect 14252 22133 14258 22167
rect 14292 22133 14298 22167
rect 14252 22095 14298 22133
rect 14252 22061 14258 22095
rect 14292 22061 14298 22095
rect 14252 22023 14298 22061
rect 14252 21989 14258 22023
rect 14292 21989 14298 22023
rect 14252 21951 14298 21989
rect 14252 21917 14258 21951
rect 14292 21917 14298 21951
rect 14252 21879 14298 21917
rect 14252 21845 14258 21879
rect 14292 21845 14298 21879
rect 14252 21807 14298 21845
rect 14252 21773 14258 21807
rect 14292 21773 14298 21807
rect 14252 21735 14298 21773
rect 14252 21701 14258 21735
rect 14292 21701 14298 21735
rect 14252 21663 14298 21701
rect 14252 21629 14258 21663
rect 14292 21629 14298 21663
rect 14252 21591 14298 21629
rect 14252 21557 14258 21591
rect 14292 21557 14298 21591
rect 14252 21519 14298 21557
rect 14252 21485 14258 21519
rect 14292 21485 14298 21519
rect 14252 21447 14298 21485
rect 14252 21413 14258 21447
rect 14292 21413 14298 21447
rect 14252 21375 14298 21413
rect 14252 21341 14258 21375
rect 14292 21341 14298 21375
rect 14252 21303 14298 21341
rect 14196 21269 14211 21271
rect 14141 21237 14211 21269
rect 14141 21185 14150 21237
rect 14202 21185 14211 21237
rect 14141 21151 14211 21185
rect 14252 21269 14258 21303
rect 14292 21269 14298 21303
rect 14348 22997 14354 23031
rect 14388 22997 14394 23031
rect 14348 22959 14394 22997
rect 14348 22925 14354 22959
rect 14388 22925 14394 22959
rect 14348 22887 14394 22925
rect 14348 22853 14354 22887
rect 14388 22853 14394 22887
rect 14348 22815 14394 22853
rect 14348 22781 14354 22815
rect 14388 22781 14394 22815
rect 14348 22743 14394 22781
rect 14348 22709 14354 22743
rect 14388 22709 14394 22743
rect 14348 22671 14394 22709
rect 14348 22637 14354 22671
rect 14388 22637 14394 22671
rect 14348 22599 14394 22637
rect 14348 22565 14354 22599
rect 14388 22565 14394 22599
rect 14348 22527 14394 22565
rect 14348 22493 14354 22527
rect 14388 22493 14394 22527
rect 14348 22455 14394 22493
rect 14348 22421 14354 22455
rect 14388 22421 14394 22455
rect 14348 22383 14394 22421
rect 14348 22349 14354 22383
rect 14388 22349 14394 22383
rect 14348 22311 14394 22349
rect 14348 22277 14354 22311
rect 14388 22277 14394 22311
rect 14348 22239 14394 22277
rect 14348 22205 14354 22239
rect 14388 22205 14394 22239
rect 14348 22167 14394 22205
rect 14348 22133 14354 22167
rect 14388 22133 14394 22167
rect 14348 22095 14394 22133
rect 14348 22061 14354 22095
rect 14388 22061 14394 22095
rect 14348 22023 14394 22061
rect 14348 21989 14354 22023
rect 14388 21989 14394 22023
rect 14348 21951 14394 21989
rect 14348 21917 14354 21951
rect 14388 21917 14394 21951
rect 14348 21879 14394 21917
rect 14348 21845 14354 21879
rect 14388 21845 14394 21879
rect 14348 21807 14394 21845
rect 14348 21773 14354 21807
rect 14388 21773 14394 21807
rect 14348 21735 14394 21773
rect 14348 21701 14354 21735
rect 14388 21701 14394 21735
rect 14348 21663 14394 21701
rect 14348 21629 14354 21663
rect 14388 21629 14394 21663
rect 14348 21591 14394 21629
rect 14348 21557 14354 21591
rect 14388 21557 14394 21591
rect 14348 21519 14394 21557
rect 14348 21485 14354 21519
rect 14388 21485 14394 21519
rect 14348 21447 14394 21485
rect 14348 21413 14354 21447
rect 14388 21413 14394 21447
rect 14348 21375 14394 21413
rect 14348 21341 14354 21375
rect 14388 21341 14394 21375
rect 14348 21303 14394 21341
rect 14348 21271 14354 21303
rect 14252 21231 14298 21269
rect 14252 21197 14258 21231
rect 14292 21197 14298 21231
rect 14156 21150 14202 21151
rect 14252 21150 14298 21197
rect 14331 21269 14354 21271
rect 14388 21271 14394 21303
rect 14444 22997 14450 23031
rect 14484 22997 14490 23031
rect 14444 22959 14490 22997
rect 14444 22925 14450 22959
rect 14484 22925 14490 22959
rect 14444 22887 14490 22925
rect 14444 22853 14450 22887
rect 14484 22853 14490 22887
rect 14444 22815 14490 22853
rect 14444 22781 14450 22815
rect 14484 22781 14490 22815
rect 14444 22743 14490 22781
rect 14444 22709 14450 22743
rect 14484 22709 14490 22743
rect 14444 22671 14490 22709
rect 14444 22637 14450 22671
rect 14484 22637 14490 22671
rect 14444 22599 14490 22637
rect 14444 22565 14450 22599
rect 14484 22565 14490 22599
rect 14444 22527 14490 22565
rect 14444 22493 14450 22527
rect 14484 22493 14490 22527
rect 14444 22455 14490 22493
rect 14444 22421 14450 22455
rect 14484 22421 14490 22455
rect 14444 22383 14490 22421
rect 14444 22349 14450 22383
rect 14484 22349 14490 22383
rect 14444 22311 14490 22349
rect 14444 22277 14450 22311
rect 14484 22277 14490 22311
rect 14444 22239 14490 22277
rect 14444 22205 14450 22239
rect 14484 22205 14490 22239
rect 14444 22167 14490 22205
rect 14444 22133 14450 22167
rect 14484 22133 14490 22167
rect 14444 22095 14490 22133
rect 14444 22061 14450 22095
rect 14484 22061 14490 22095
rect 14444 22023 14490 22061
rect 14444 21989 14450 22023
rect 14484 21989 14490 22023
rect 14444 21951 14490 21989
rect 14444 21917 14450 21951
rect 14484 21917 14490 21951
rect 14444 21879 14490 21917
rect 14444 21845 14450 21879
rect 14484 21845 14490 21879
rect 14444 21807 14490 21845
rect 14444 21773 14450 21807
rect 14484 21773 14490 21807
rect 14444 21735 14490 21773
rect 14444 21701 14450 21735
rect 14484 21701 14490 21735
rect 14444 21663 14490 21701
rect 14444 21629 14450 21663
rect 14484 21629 14490 21663
rect 14444 21591 14490 21629
rect 14444 21557 14450 21591
rect 14484 21557 14490 21591
rect 14444 21519 14490 21557
rect 14444 21485 14450 21519
rect 14484 21485 14490 21519
rect 14444 21447 14490 21485
rect 14444 21413 14450 21447
rect 14484 21413 14490 21447
rect 14444 21375 14490 21413
rect 14444 21341 14450 21375
rect 14484 21341 14490 21375
rect 14444 21303 14490 21341
rect 14388 21269 14401 21271
rect 14331 21237 14401 21269
rect 14331 21185 14340 21237
rect 14392 21185 14401 21237
rect 14331 21151 14401 21185
rect 14444 21269 14450 21303
rect 14484 21269 14490 21303
rect 14540 22997 14546 23031
rect 14580 22997 14586 23031
rect 14540 22959 14586 22997
rect 14540 22925 14546 22959
rect 14580 22925 14586 22959
rect 14540 22887 14586 22925
rect 14540 22853 14546 22887
rect 14580 22853 14586 22887
rect 14540 22815 14586 22853
rect 14540 22781 14546 22815
rect 14580 22781 14586 22815
rect 14540 22743 14586 22781
rect 14540 22709 14546 22743
rect 14580 22709 14586 22743
rect 14540 22671 14586 22709
rect 14540 22637 14546 22671
rect 14580 22637 14586 22671
rect 14540 22599 14586 22637
rect 14540 22565 14546 22599
rect 14580 22565 14586 22599
rect 14540 22527 14586 22565
rect 14540 22493 14546 22527
rect 14580 22493 14586 22527
rect 14540 22455 14586 22493
rect 14540 22421 14546 22455
rect 14580 22421 14586 22455
rect 14540 22383 14586 22421
rect 14540 22349 14546 22383
rect 14580 22349 14586 22383
rect 14540 22311 14586 22349
rect 14540 22277 14546 22311
rect 14580 22277 14586 22311
rect 14540 22239 14586 22277
rect 14540 22205 14546 22239
rect 14580 22205 14586 22239
rect 14540 22167 14586 22205
rect 14540 22133 14546 22167
rect 14580 22133 14586 22167
rect 14540 22095 14586 22133
rect 14540 22061 14546 22095
rect 14580 22061 14586 22095
rect 14540 22023 14586 22061
rect 14540 21989 14546 22023
rect 14580 21989 14586 22023
rect 14540 21951 14586 21989
rect 14540 21917 14546 21951
rect 14580 21917 14586 21951
rect 14540 21879 14586 21917
rect 14540 21845 14546 21879
rect 14580 21845 14586 21879
rect 14540 21807 14586 21845
rect 14540 21773 14546 21807
rect 14580 21773 14586 21807
rect 14540 21735 14586 21773
rect 14540 21701 14546 21735
rect 14580 21701 14586 21735
rect 14540 21663 14586 21701
rect 14540 21629 14546 21663
rect 14580 21629 14586 21663
rect 14540 21591 14586 21629
rect 14540 21557 14546 21591
rect 14580 21557 14586 21591
rect 14540 21519 14586 21557
rect 14540 21485 14546 21519
rect 14580 21485 14586 21519
rect 14540 21447 14586 21485
rect 14540 21413 14546 21447
rect 14580 21413 14586 21447
rect 14540 21375 14586 21413
rect 14540 21341 14546 21375
rect 14580 21341 14586 21375
rect 14540 21303 14586 21341
rect 14540 21271 14546 21303
rect 14444 21231 14490 21269
rect 14444 21197 14450 21231
rect 14484 21197 14490 21231
rect 14348 21150 14394 21151
rect 14444 21150 14490 21197
rect 14521 21269 14546 21271
rect 14580 21271 14586 21303
rect 14636 22997 14642 23031
rect 14676 22997 14682 23031
rect 14636 22959 14682 22997
rect 14636 22925 14642 22959
rect 14676 22925 14682 22959
rect 14636 22887 14682 22925
rect 14636 22853 14642 22887
rect 14676 22853 14682 22887
rect 14636 22815 14682 22853
rect 14636 22781 14642 22815
rect 14676 22781 14682 22815
rect 14636 22743 14682 22781
rect 14636 22709 14642 22743
rect 14676 22709 14682 22743
rect 14636 22671 14682 22709
rect 14636 22637 14642 22671
rect 14676 22637 14682 22671
rect 14636 22599 14682 22637
rect 14636 22565 14642 22599
rect 14676 22565 14682 22599
rect 14636 22527 14682 22565
rect 14636 22493 14642 22527
rect 14676 22493 14682 22527
rect 14636 22455 14682 22493
rect 14636 22421 14642 22455
rect 14676 22421 14682 22455
rect 14636 22383 14682 22421
rect 14636 22349 14642 22383
rect 14676 22349 14682 22383
rect 14636 22311 14682 22349
rect 14636 22277 14642 22311
rect 14676 22277 14682 22311
rect 14636 22239 14682 22277
rect 14636 22205 14642 22239
rect 14676 22205 14682 22239
rect 14636 22167 14682 22205
rect 14636 22133 14642 22167
rect 14676 22133 14682 22167
rect 14636 22095 14682 22133
rect 14636 22061 14642 22095
rect 14676 22061 14682 22095
rect 14636 22023 14682 22061
rect 14636 21989 14642 22023
rect 14676 21989 14682 22023
rect 14636 21951 14682 21989
rect 14636 21917 14642 21951
rect 14676 21917 14682 21951
rect 14636 21879 14682 21917
rect 14636 21845 14642 21879
rect 14676 21845 14682 21879
rect 14636 21807 14682 21845
rect 14636 21773 14642 21807
rect 14676 21773 14682 21807
rect 14636 21735 14682 21773
rect 14636 21701 14642 21735
rect 14676 21701 14682 21735
rect 14636 21663 14682 21701
rect 14636 21629 14642 21663
rect 14676 21629 14682 21663
rect 14636 21591 14682 21629
rect 14636 21557 14642 21591
rect 14676 21557 14682 21591
rect 14636 21519 14682 21557
rect 14636 21485 14642 21519
rect 14676 21485 14682 21519
rect 14636 21447 14682 21485
rect 14636 21413 14642 21447
rect 14676 21413 14682 21447
rect 14636 21375 14682 21413
rect 14636 21341 14642 21375
rect 14676 21341 14682 21375
rect 14636 21303 14682 21341
rect 14580 21269 14591 21271
rect 14521 21237 14591 21269
rect 14521 21185 14530 21237
rect 14582 21185 14591 21237
rect 14521 21151 14591 21185
rect 14636 21269 14642 21303
rect 14676 21269 14682 21303
rect 14732 22997 14738 23031
rect 14772 22997 14778 23031
rect 14810 23116 14920 23160
rect 14810 23064 14839 23116
rect 14891 23064 14920 23116
rect 14810 23020 14920 23064
rect 15260 23138 15420 23176
rect 15260 23104 15324 23138
rect 15358 23104 15420 23138
rect 15260 23066 15420 23104
rect 15260 23032 15324 23066
rect 15358 23032 15420 23066
rect 14732 22959 14778 22997
rect 14732 22925 14738 22959
rect 14772 22925 14778 22959
rect 14732 22887 14778 22925
rect 14732 22853 14738 22887
rect 14772 22853 14778 22887
rect 14732 22815 14778 22853
rect 14732 22781 14738 22815
rect 14772 22781 14778 22815
rect 14732 22743 14778 22781
rect 15260 22994 15420 23032
rect 15260 22960 15324 22994
rect 15358 22960 15420 22994
rect 15260 22922 15420 22960
rect 15260 22888 15324 22922
rect 15358 22888 15420 22922
rect 15260 22850 15420 22888
rect 15260 22816 15324 22850
rect 15358 22816 15420 22850
rect 15260 22760 15420 22816
rect 15824 23142 15870 23189
rect 15824 23108 15830 23142
rect 15864 23108 15870 23142
rect 15824 23070 15870 23108
rect 15901 23157 15971 23191
rect 15901 23105 15910 23157
rect 15962 23105 15971 23157
rect 15901 23071 15971 23105
rect 16016 23142 16062 23189
rect 16016 23108 16022 23142
rect 16056 23108 16062 23142
rect 15824 23036 15830 23070
rect 15864 23036 15870 23070
rect 15824 22998 15870 23036
rect 15824 22964 15830 22998
rect 15864 22964 15870 22998
rect 15824 22926 15870 22964
rect 15824 22892 15830 22926
rect 15864 22892 15870 22926
rect 15824 22854 15870 22892
rect 15824 22820 15830 22854
rect 15864 22820 15870 22854
rect 15824 22782 15870 22820
rect 14732 22709 14738 22743
rect 14772 22709 14778 22743
rect 14732 22671 14778 22709
rect 14732 22637 14738 22671
rect 14772 22637 14778 22671
rect 14732 22599 14778 22637
rect 14732 22565 14738 22599
rect 14772 22565 14778 22599
rect 14732 22527 14778 22565
rect 14732 22493 14738 22527
rect 14772 22493 14778 22527
rect 14732 22455 14778 22493
rect 14732 22421 14738 22455
rect 14772 22421 14778 22455
rect 14732 22383 14778 22421
rect 14732 22349 14738 22383
rect 14772 22349 14778 22383
rect 14732 22311 14778 22349
rect 14732 22277 14738 22311
rect 14772 22277 14778 22311
rect 14732 22239 14778 22277
rect 14732 22205 14738 22239
rect 14772 22205 14778 22239
rect 14732 22167 14778 22205
rect 14732 22133 14738 22167
rect 14772 22133 14778 22167
rect 14732 22095 14778 22133
rect 14732 22061 14738 22095
rect 14772 22061 14778 22095
rect 14732 22023 14778 22061
rect 14732 21989 14738 22023
rect 14772 21989 14778 22023
rect 14732 21951 14778 21989
rect 14732 21917 14738 21951
rect 14772 21917 14778 21951
rect 14732 21879 14778 21917
rect 14732 21845 14738 21879
rect 14772 21845 14778 21879
rect 14732 21807 14778 21845
rect 14732 21773 14738 21807
rect 14772 21773 14778 21807
rect 14732 21735 14778 21773
rect 14732 21701 14738 21735
rect 14772 21701 14778 21735
rect 14732 21663 14778 21701
rect 14732 21629 14738 21663
rect 14772 21629 14778 21663
rect 14732 21591 14778 21629
rect 14732 21557 14738 21591
rect 14772 21557 14778 21591
rect 14732 21519 14778 21557
rect 15824 22748 15830 22782
rect 15864 22748 15870 22782
rect 15824 22710 15870 22748
rect 15824 22676 15830 22710
rect 15864 22676 15870 22710
rect 15824 22638 15870 22676
rect 15824 22604 15830 22638
rect 15864 22604 15870 22638
rect 15824 22566 15870 22604
rect 15824 22532 15830 22566
rect 15864 22532 15870 22566
rect 15824 22494 15870 22532
rect 15824 22460 15830 22494
rect 15864 22460 15870 22494
rect 15824 22422 15870 22460
rect 15824 22388 15830 22422
rect 15864 22388 15870 22422
rect 15824 22350 15870 22388
rect 15824 22316 15830 22350
rect 15864 22316 15870 22350
rect 15824 22278 15870 22316
rect 15824 22244 15830 22278
rect 15864 22244 15870 22278
rect 15824 22206 15870 22244
rect 15824 22172 15830 22206
rect 15864 22172 15870 22206
rect 15824 22134 15870 22172
rect 15824 22100 15830 22134
rect 15864 22100 15870 22134
rect 15824 22062 15870 22100
rect 15824 22028 15830 22062
rect 15864 22028 15870 22062
rect 15824 21990 15870 22028
rect 15824 21956 15830 21990
rect 15864 21956 15870 21990
rect 15824 21918 15870 21956
rect 15824 21884 15830 21918
rect 15864 21884 15870 21918
rect 15824 21846 15870 21884
rect 15824 21812 15830 21846
rect 15864 21812 15870 21846
rect 15824 21774 15870 21812
rect 15824 21740 15830 21774
rect 15864 21740 15870 21774
rect 15824 21702 15870 21740
rect 15824 21668 15830 21702
rect 15864 21668 15870 21702
rect 15824 21630 15870 21668
rect 15824 21596 15830 21630
rect 15864 21596 15870 21630
rect 15824 21558 15870 21596
rect 14732 21485 14738 21519
rect 14772 21485 14778 21519
rect 14732 21447 14778 21485
rect 14732 21413 14738 21447
rect 14772 21413 14778 21447
rect 14732 21375 14778 21413
rect 14732 21341 14738 21375
rect 14772 21341 14778 21375
rect 14732 21303 14778 21341
rect 14732 21271 14738 21303
rect 14636 21231 14682 21269
rect 14636 21197 14642 21231
rect 14676 21197 14682 21231
rect 14540 21150 14586 21151
rect 14636 21150 14682 21197
rect 14721 21269 14738 21271
rect 14772 21271 14778 21303
rect 15316 21539 15366 21553
rect 15316 21505 15324 21539
rect 15358 21505 15366 21539
rect 15316 21467 15366 21505
rect 15316 21433 15324 21467
rect 15358 21433 15366 21467
rect 15316 21395 15366 21433
rect 15316 21361 15324 21395
rect 15358 21361 15366 21395
rect 15316 21323 15366 21361
rect 15316 21290 15324 21323
rect 15290 21289 15324 21290
rect 15358 21290 15366 21323
rect 15824 21524 15830 21558
rect 15864 21524 15870 21558
rect 15824 21486 15870 21524
rect 15824 21452 15830 21486
rect 15864 21452 15870 21486
rect 15824 21414 15870 21452
rect 15824 21380 15830 21414
rect 15864 21380 15870 21414
rect 15824 21342 15870 21380
rect 15824 21311 15830 21342
rect 15801 21308 15830 21311
rect 15864 21311 15870 21342
rect 15920 23070 15966 23071
rect 15920 23036 15926 23070
rect 15960 23036 15966 23070
rect 15920 22998 15966 23036
rect 15920 22964 15926 22998
rect 15960 22964 15966 22998
rect 15920 22926 15966 22964
rect 15920 22892 15926 22926
rect 15960 22892 15966 22926
rect 15920 22854 15966 22892
rect 15920 22820 15926 22854
rect 15960 22820 15966 22854
rect 15920 22782 15966 22820
rect 15920 22748 15926 22782
rect 15960 22748 15966 22782
rect 15920 22710 15966 22748
rect 15920 22676 15926 22710
rect 15960 22676 15966 22710
rect 15920 22638 15966 22676
rect 15920 22604 15926 22638
rect 15960 22604 15966 22638
rect 15920 22566 15966 22604
rect 15920 22532 15926 22566
rect 15960 22532 15966 22566
rect 15920 22494 15966 22532
rect 15920 22460 15926 22494
rect 15960 22460 15966 22494
rect 15920 22422 15966 22460
rect 15920 22388 15926 22422
rect 15960 22388 15966 22422
rect 15920 22350 15966 22388
rect 15920 22316 15926 22350
rect 15960 22316 15966 22350
rect 15920 22278 15966 22316
rect 15920 22244 15926 22278
rect 15960 22244 15966 22278
rect 15920 22206 15966 22244
rect 15920 22172 15926 22206
rect 15960 22172 15966 22206
rect 15920 22134 15966 22172
rect 15920 22100 15926 22134
rect 15960 22100 15966 22134
rect 15920 22062 15966 22100
rect 15920 22028 15926 22062
rect 15960 22028 15966 22062
rect 15920 21990 15966 22028
rect 15920 21956 15926 21990
rect 15960 21956 15966 21990
rect 15920 21918 15966 21956
rect 15920 21884 15926 21918
rect 15960 21884 15966 21918
rect 15920 21846 15966 21884
rect 15920 21812 15926 21846
rect 15960 21812 15966 21846
rect 15920 21774 15966 21812
rect 15920 21740 15926 21774
rect 15960 21740 15966 21774
rect 15920 21702 15966 21740
rect 15920 21668 15926 21702
rect 15960 21668 15966 21702
rect 15920 21630 15966 21668
rect 15920 21596 15926 21630
rect 15960 21596 15966 21630
rect 15920 21558 15966 21596
rect 15920 21524 15926 21558
rect 15960 21524 15966 21558
rect 15920 21486 15966 21524
rect 15920 21452 15926 21486
rect 15960 21452 15966 21486
rect 15920 21414 15966 21452
rect 15920 21380 15926 21414
rect 15960 21380 15966 21414
rect 15920 21342 15966 21380
rect 15864 21308 15871 21311
rect 15358 21289 15390 21290
rect 14772 21269 14791 21271
rect 14721 21237 14791 21269
rect 14721 21185 14730 21237
rect 14782 21185 14791 21237
rect 14721 21151 14791 21185
rect 15290 21251 15390 21289
rect 15290 21217 15324 21251
rect 15358 21217 15390 21251
rect 15290 21179 15390 21217
rect 15801 21277 15871 21308
rect 15801 21225 15810 21277
rect 15862 21270 15871 21277
rect 15864 21236 15871 21270
rect 15862 21225 15871 21236
rect 15801 21191 15871 21225
rect 15920 21308 15926 21342
rect 15960 21308 15966 21342
rect 16016 23070 16062 23108
rect 16091 23157 16161 23191
rect 16091 23105 16100 23157
rect 16152 23105 16161 23157
rect 16091 23071 16161 23105
rect 16656 23167 16662 23201
rect 16696 23167 16702 23201
rect 16656 23129 16702 23167
rect 16656 23095 16662 23129
rect 16696 23095 16702 23129
rect 16016 23036 16022 23070
rect 16056 23036 16062 23070
rect 16016 22998 16062 23036
rect 16016 22964 16022 22998
rect 16056 22964 16062 22998
rect 16016 22926 16062 22964
rect 16016 22892 16022 22926
rect 16056 22892 16062 22926
rect 16016 22854 16062 22892
rect 16016 22820 16022 22854
rect 16056 22820 16062 22854
rect 16016 22782 16062 22820
rect 16016 22748 16022 22782
rect 16056 22748 16062 22782
rect 16016 22710 16062 22748
rect 16016 22676 16022 22710
rect 16056 22676 16062 22710
rect 16016 22638 16062 22676
rect 16016 22604 16022 22638
rect 16056 22604 16062 22638
rect 16016 22566 16062 22604
rect 16016 22532 16022 22566
rect 16056 22532 16062 22566
rect 16016 22494 16062 22532
rect 16016 22460 16022 22494
rect 16056 22460 16062 22494
rect 16016 22422 16062 22460
rect 16016 22388 16022 22422
rect 16056 22388 16062 22422
rect 16016 22350 16062 22388
rect 16016 22316 16022 22350
rect 16056 22316 16062 22350
rect 16016 22278 16062 22316
rect 16016 22244 16022 22278
rect 16056 22244 16062 22278
rect 16016 22206 16062 22244
rect 16016 22172 16022 22206
rect 16056 22172 16062 22206
rect 16016 22134 16062 22172
rect 16016 22100 16022 22134
rect 16056 22100 16062 22134
rect 16016 22062 16062 22100
rect 16016 22028 16022 22062
rect 16056 22028 16062 22062
rect 16016 21990 16062 22028
rect 16016 21956 16022 21990
rect 16056 21956 16062 21990
rect 16016 21918 16062 21956
rect 16016 21884 16022 21918
rect 16056 21884 16062 21918
rect 16016 21846 16062 21884
rect 16016 21812 16022 21846
rect 16056 21812 16062 21846
rect 16016 21774 16062 21812
rect 16016 21740 16022 21774
rect 16056 21740 16062 21774
rect 16016 21702 16062 21740
rect 16016 21668 16022 21702
rect 16056 21668 16062 21702
rect 16016 21630 16062 21668
rect 16016 21596 16022 21630
rect 16056 21596 16062 21630
rect 16016 21558 16062 21596
rect 16016 21524 16022 21558
rect 16056 21524 16062 21558
rect 16016 21486 16062 21524
rect 16016 21452 16022 21486
rect 16056 21452 16062 21486
rect 16016 21414 16062 21452
rect 16016 21380 16022 21414
rect 16056 21380 16062 21414
rect 16016 21342 16062 21380
rect 16016 21311 16022 21342
rect 15920 21270 15966 21308
rect 15920 21236 15926 21270
rect 15960 21236 15966 21270
rect 15824 21189 15870 21191
rect 15920 21189 15966 21236
rect 16001 21308 16022 21311
rect 16056 21311 16062 21342
rect 16112 23070 16158 23071
rect 16112 23036 16118 23070
rect 16152 23036 16158 23070
rect 16112 22998 16158 23036
rect 16112 22964 16118 22998
rect 16152 22964 16158 22998
rect 16112 22926 16158 22964
rect 16112 22892 16118 22926
rect 16152 22892 16158 22926
rect 16112 22854 16158 22892
rect 16112 22820 16118 22854
rect 16152 22820 16158 22854
rect 16112 22782 16158 22820
rect 16112 22748 16118 22782
rect 16152 22748 16158 22782
rect 16112 22710 16158 22748
rect 16112 22676 16118 22710
rect 16152 22676 16158 22710
rect 16112 22638 16158 22676
rect 16112 22604 16118 22638
rect 16152 22604 16158 22638
rect 16112 22566 16158 22604
rect 16112 22532 16118 22566
rect 16152 22532 16158 22566
rect 16112 22494 16158 22532
rect 16112 22460 16118 22494
rect 16152 22460 16158 22494
rect 16112 22422 16158 22460
rect 16112 22388 16118 22422
rect 16152 22388 16158 22422
rect 16112 22350 16158 22388
rect 16112 22316 16118 22350
rect 16152 22316 16158 22350
rect 16112 22278 16158 22316
rect 16112 22244 16118 22278
rect 16152 22244 16158 22278
rect 16112 22206 16158 22244
rect 16112 22172 16118 22206
rect 16152 22172 16158 22206
rect 16112 22134 16158 22172
rect 16656 23057 16702 23095
rect 16656 23023 16662 23057
rect 16696 23023 16702 23057
rect 16656 22985 16702 23023
rect 16656 22951 16662 22985
rect 16696 22951 16702 22985
rect 16656 22913 16702 22951
rect 16656 22879 16662 22913
rect 16696 22879 16702 22913
rect 16656 22841 16702 22879
rect 16656 22807 16662 22841
rect 16696 22807 16702 22841
rect 16656 22769 16702 22807
rect 16656 22735 16662 22769
rect 16696 22735 16702 22769
rect 16656 22697 16702 22735
rect 16656 22663 16662 22697
rect 16696 22663 16702 22697
rect 16656 22625 16702 22663
rect 16656 22591 16662 22625
rect 16696 22591 16702 22625
rect 16656 22553 16702 22591
rect 16656 22519 16662 22553
rect 16696 22519 16702 22553
rect 16656 22481 16702 22519
rect 16656 22447 16662 22481
rect 16696 22447 16702 22481
rect 16656 22409 16702 22447
rect 16656 22375 16662 22409
rect 16696 22375 16702 22409
rect 16656 22337 16702 22375
rect 16656 22303 16662 22337
rect 16696 22303 16702 22337
rect 16656 22265 16702 22303
rect 16656 22231 16662 22265
rect 16696 22231 16702 22265
rect 16656 22193 16702 22231
rect 16656 22170 16662 22193
rect 16112 22100 16118 22134
rect 16152 22100 16158 22134
rect 16112 22062 16158 22100
rect 16112 22028 16118 22062
rect 16152 22028 16158 22062
rect 16651 22159 16662 22170
rect 16696 22170 16702 22193
rect 16752 23887 16758 23911
rect 16792 23911 16813 23921
rect 16848 23993 16894 24040
rect 16848 23959 16854 23993
rect 16888 23959 16894 23993
rect 16848 23921 16894 23959
rect 16792 23887 16798 23911
rect 16752 23849 16798 23887
rect 16752 23815 16758 23849
rect 16792 23815 16798 23849
rect 16752 23777 16798 23815
rect 16752 23743 16758 23777
rect 16792 23743 16798 23777
rect 16752 23705 16798 23743
rect 16752 23671 16758 23705
rect 16792 23671 16798 23705
rect 16752 23633 16798 23671
rect 16752 23599 16758 23633
rect 16792 23599 16798 23633
rect 16752 23561 16798 23599
rect 16752 23527 16758 23561
rect 16792 23527 16798 23561
rect 16752 23489 16798 23527
rect 16752 23455 16758 23489
rect 16792 23455 16798 23489
rect 16752 23417 16798 23455
rect 16752 23383 16758 23417
rect 16792 23383 16798 23417
rect 16752 23345 16798 23383
rect 16752 23311 16758 23345
rect 16792 23311 16798 23345
rect 16752 23273 16798 23311
rect 16752 23239 16758 23273
rect 16792 23239 16798 23273
rect 16752 23201 16798 23239
rect 16752 23167 16758 23201
rect 16792 23167 16798 23201
rect 16752 23129 16798 23167
rect 16752 23095 16758 23129
rect 16792 23095 16798 23129
rect 16752 23057 16798 23095
rect 16752 23023 16758 23057
rect 16792 23023 16798 23057
rect 16752 22985 16798 23023
rect 16752 22951 16758 22985
rect 16792 22951 16798 22985
rect 16752 22913 16798 22951
rect 16752 22879 16758 22913
rect 16792 22879 16798 22913
rect 16752 22841 16798 22879
rect 16752 22807 16758 22841
rect 16792 22807 16798 22841
rect 16752 22769 16798 22807
rect 16752 22735 16758 22769
rect 16792 22735 16798 22769
rect 16752 22697 16798 22735
rect 16752 22663 16758 22697
rect 16792 22663 16798 22697
rect 16752 22625 16798 22663
rect 16752 22591 16758 22625
rect 16792 22591 16798 22625
rect 16752 22553 16798 22591
rect 16752 22519 16758 22553
rect 16792 22519 16798 22553
rect 16752 22481 16798 22519
rect 16752 22447 16758 22481
rect 16792 22447 16798 22481
rect 16752 22409 16798 22447
rect 16752 22375 16758 22409
rect 16792 22375 16798 22409
rect 16752 22337 16798 22375
rect 16752 22303 16758 22337
rect 16792 22303 16798 22337
rect 16752 22265 16798 22303
rect 16752 22231 16758 22265
rect 16792 22231 16798 22265
rect 16752 22193 16798 22231
rect 16696 22159 16721 22170
rect 16651 22130 16721 22159
rect 16651 22078 16658 22130
rect 16710 22078 16721 22130
rect 16651 22040 16721 22078
rect 16752 22159 16758 22193
rect 16792 22159 16798 22193
rect 16848 23887 16854 23921
rect 16888 23887 16894 23921
rect 16933 24001 17003 24041
rect 16933 23949 16940 24001
rect 16992 23949 17003 24001
rect 16933 23921 17003 23949
rect 16933 23911 16950 23921
rect 16848 23849 16894 23887
rect 16848 23815 16854 23849
rect 16888 23815 16894 23849
rect 16848 23777 16894 23815
rect 16848 23743 16854 23777
rect 16888 23743 16894 23777
rect 16848 23705 16894 23743
rect 16848 23671 16854 23705
rect 16888 23671 16894 23705
rect 16848 23633 16894 23671
rect 16848 23599 16854 23633
rect 16888 23599 16894 23633
rect 16848 23561 16894 23599
rect 16848 23527 16854 23561
rect 16888 23527 16894 23561
rect 16848 23489 16894 23527
rect 16848 23455 16854 23489
rect 16888 23455 16894 23489
rect 16848 23417 16894 23455
rect 16848 23383 16854 23417
rect 16888 23383 16894 23417
rect 16848 23345 16894 23383
rect 16848 23311 16854 23345
rect 16888 23311 16894 23345
rect 16848 23273 16894 23311
rect 16848 23239 16854 23273
rect 16888 23239 16894 23273
rect 16848 23201 16894 23239
rect 16848 23167 16854 23201
rect 16888 23167 16894 23201
rect 16848 23129 16894 23167
rect 16848 23095 16854 23129
rect 16888 23095 16894 23129
rect 16848 23057 16894 23095
rect 16848 23023 16854 23057
rect 16888 23023 16894 23057
rect 16848 22985 16894 23023
rect 16848 22951 16854 22985
rect 16888 22951 16894 22985
rect 16848 22913 16894 22951
rect 16848 22879 16854 22913
rect 16888 22879 16894 22913
rect 16848 22841 16894 22879
rect 16848 22807 16854 22841
rect 16888 22807 16894 22841
rect 16848 22769 16894 22807
rect 16848 22735 16854 22769
rect 16888 22735 16894 22769
rect 16848 22697 16894 22735
rect 16848 22663 16854 22697
rect 16888 22663 16894 22697
rect 16848 22625 16894 22663
rect 16848 22591 16854 22625
rect 16888 22591 16894 22625
rect 16848 22553 16894 22591
rect 16848 22519 16854 22553
rect 16888 22519 16894 22553
rect 16848 22481 16894 22519
rect 16848 22447 16854 22481
rect 16888 22447 16894 22481
rect 16848 22409 16894 22447
rect 16848 22375 16854 22409
rect 16888 22375 16894 22409
rect 16848 22337 16894 22375
rect 16848 22303 16854 22337
rect 16888 22303 16894 22337
rect 16848 22265 16894 22303
rect 16848 22231 16854 22265
rect 16888 22231 16894 22265
rect 16848 22193 16894 22231
rect 16848 22170 16854 22193
rect 16752 22121 16798 22159
rect 16752 22087 16758 22121
rect 16792 22087 16798 22121
rect 16752 22040 16798 22087
rect 16832 22159 16854 22170
rect 16888 22170 16894 22193
rect 16944 23887 16950 23911
rect 16984 23911 17003 23921
rect 17040 23993 17086 24040
rect 17040 23959 17046 23993
rect 17080 23959 17086 23993
rect 17040 23921 17086 23959
rect 16984 23887 16990 23911
rect 16944 23849 16990 23887
rect 16944 23815 16950 23849
rect 16984 23815 16990 23849
rect 16944 23777 16990 23815
rect 16944 23743 16950 23777
rect 16984 23743 16990 23777
rect 16944 23705 16990 23743
rect 16944 23671 16950 23705
rect 16984 23671 16990 23705
rect 16944 23633 16990 23671
rect 16944 23599 16950 23633
rect 16984 23599 16990 23633
rect 16944 23561 16990 23599
rect 16944 23527 16950 23561
rect 16984 23527 16990 23561
rect 16944 23489 16990 23527
rect 16944 23455 16950 23489
rect 16984 23455 16990 23489
rect 16944 23417 16990 23455
rect 16944 23383 16950 23417
rect 16984 23383 16990 23417
rect 16944 23345 16990 23383
rect 16944 23311 16950 23345
rect 16984 23311 16990 23345
rect 16944 23273 16990 23311
rect 16944 23239 16950 23273
rect 16984 23239 16990 23273
rect 16944 23201 16990 23239
rect 16944 23167 16950 23201
rect 16984 23167 16990 23201
rect 16944 23129 16990 23167
rect 16944 23095 16950 23129
rect 16984 23095 16990 23129
rect 16944 23057 16990 23095
rect 16944 23023 16950 23057
rect 16984 23023 16990 23057
rect 16944 22985 16990 23023
rect 16944 22951 16950 22985
rect 16984 22951 16990 22985
rect 16944 22913 16990 22951
rect 16944 22879 16950 22913
rect 16984 22879 16990 22913
rect 16944 22841 16990 22879
rect 16944 22807 16950 22841
rect 16984 22807 16990 22841
rect 16944 22769 16990 22807
rect 16944 22735 16950 22769
rect 16984 22735 16990 22769
rect 16944 22697 16990 22735
rect 16944 22663 16950 22697
rect 16984 22663 16990 22697
rect 16944 22625 16990 22663
rect 16944 22591 16950 22625
rect 16984 22591 16990 22625
rect 16944 22553 16990 22591
rect 16944 22519 16950 22553
rect 16984 22519 16990 22553
rect 16944 22481 16990 22519
rect 16944 22447 16950 22481
rect 16984 22447 16990 22481
rect 16944 22409 16990 22447
rect 16944 22375 16950 22409
rect 16984 22375 16990 22409
rect 16944 22337 16990 22375
rect 16944 22303 16950 22337
rect 16984 22303 16990 22337
rect 16944 22265 16990 22303
rect 16944 22231 16950 22265
rect 16984 22231 16990 22265
rect 16944 22193 16990 22231
rect 16888 22159 16902 22170
rect 16832 22130 16902 22159
rect 16832 22078 16839 22130
rect 16891 22078 16902 22130
rect 16832 22040 16902 22078
rect 16944 22159 16950 22193
rect 16984 22159 16990 22193
rect 17040 23887 17046 23921
rect 17080 23887 17086 23921
rect 17123 24001 17193 24041
rect 17123 23949 17130 24001
rect 17182 23949 17193 24001
rect 17123 23921 17193 23949
rect 17123 23911 17142 23921
rect 17040 23849 17086 23887
rect 17040 23815 17046 23849
rect 17080 23815 17086 23849
rect 17040 23777 17086 23815
rect 17040 23743 17046 23777
rect 17080 23743 17086 23777
rect 17040 23705 17086 23743
rect 17040 23671 17046 23705
rect 17080 23671 17086 23705
rect 17040 23633 17086 23671
rect 17040 23599 17046 23633
rect 17080 23599 17086 23633
rect 17040 23561 17086 23599
rect 17040 23527 17046 23561
rect 17080 23527 17086 23561
rect 17040 23489 17086 23527
rect 17040 23455 17046 23489
rect 17080 23455 17086 23489
rect 17040 23417 17086 23455
rect 17040 23383 17046 23417
rect 17080 23383 17086 23417
rect 17040 23345 17086 23383
rect 17040 23311 17046 23345
rect 17080 23311 17086 23345
rect 17040 23273 17086 23311
rect 17040 23239 17046 23273
rect 17080 23239 17086 23273
rect 17040 23201 17086 23239
rect 17040 23167 17046 23201
rect 17080 23167 17086 23201
rect 17040 23129 17086 23167
rect 17040 23095 17046 23129
rect 17080 23095 17086 23129
rect 17040 23057 17086 23095
rect 17040 23023 17046 23057
rect 17080 23023 17086 23057
rect 17040 22985 17086 23023
rect 17040 22951 17046 22985
rect 17080 22951 17086 22985
rect 17040 22913 17086 22951
rect 17040 22879 17046 22913
rect 17080 22879 17086 22913
rect 17040 22841 17086 22879
rect 17040 22807 17046 22841
rect 17080 22807 17086 22841
rect 17040 22769 17086 22807
rect 17040 22735 17046 22769
rect 17080 22735 17086 22769
rect 17040 22697 17086 22735
rect 17040 22663 17046 22697
rect 17080 22663 17086 22697
rect 17040 22625 17086 22663
rect 17040 22591 17046 22625
rect 17080 22591 17086 22625
rect 17040 22553 17086 22591
rect 17040 22519 17046 22553
rect 17080 22519 17086 22553
rect 17040 22481 17086 22519
rect 17040 22447 17046 22481
rect 17080 22447 17086 22481
rect 17040 22409 17086 22447
rect 17040 22375 17046 22409
rect 17080 22375 17086 22409
rect 17040 22337 17086 22375
rect 17040 22303 17046 22337
rect 17080 22303 17086 22337
rect 17040 22265 17086 22303
rect 17040 22231 17046 22265
rect 17080 22231 17086 22265
rect 17040 22193 17086 22231
rect 17040 22170 17046 22193
rect 16944 22121 16990 22159
rect 16944 22087 16950 22121
rect 16984 22087 16990 22121
rect 16944 22040 16990 22087
rect 17022 22159 17046 22170
rect 17080 22170 17086 22193
rect 17136 23887 17142 23911
rect 17176 23911 17193 23921
rect 17232 23993 17278 24040
rect 17232 23959 17238 23993
rect 17272 23959 17278 23993
rect 17232 23921 17278 23959
rect 17176 23887 17182 23911
rect 17136 23849 17182 23887
rect 17136 23815 17142 23849
rect 17176 23815 17182 23849
rect 17136 23777 17182 23815
rect 17136 23743 17142 23777
rect 17176 23743 17182 23777
rect 17136 23705 17182 23743
rect 17136 23671 17142 23705
rect 17176 23671 17182 23705
rect 17136 23633 17182 23671
rect 17136 23599 17142 23633
rect 17176 23599 17182 23633
rect 17136 23561 17182 23599
rect 17136 23527 17142 23561
rect 17176 23527 17182 23561
rect 17136 23489 17182 23527
rect 17136 23455 17142 23489
rect 17176 23455 17182 23489
rect 17136 23417 17182 23455
rect 17136 23383 17142 23417
rect 17176 23383 17182 23417
rect 17136 23345 17182 23383
rect 17136 23311 17142 23345
rect 17176 23311 17182 23345
rect 17136 23273 17182 23311
rect 17136 23239 17142 23273
rect 17176 23239 17182 23273
rect 17136 23201 17182 23239
rect 17136 23167 17142 23201
rect 17176 23167 17182 23201
rect 17136 23129 17182 23167
rect 17136 23095 17142 23129
rect 17176 23095 17182 23129
rect 17136 23057 17182 23095
rect 17136 23023 17142 23057
rect 17176 23023 17182 23057
rect 17136 22985 17182 23023
rect 17136 22951 17142 22985
rect 17176 22951 17182 22985
rect 17136 22913 17182 22951
rect 17136 22879 17142 22913
rect 17176 22879 17182 22913
rect 17136 22841 17182 22879
rect 17136 22807 17142 22841
rect 17176 22807 17182 22841
rect 17136 22769 17182 22807
rect 17136 22735 17142 22769
rect 17176 22735 17182 22769
rect 17136 22697 17182 22735
rect 17136 22663 17142 22697
rect 17176 22663 17182 22697
rect 17136 22625 17182 22663
rect 17136 22591 17142 22625
rect 17176 22591 17182 22625
rect 17136 22553 17182 22591
rect 17136 22519 17142 22553
rect 17176 22519 17182 22553
rect 17136 22481 17182 22519
rect 17136 22447 17142 22481
rect 17176 22447 17182 22481
rect 17136 22409 17182 22447
rect 17136 22375 17142 22409
rect 17176 22375 17182 22409
rect 17136 22337 17182 22375
rect 17136 22303 17142 22337
rect 17176 22303 17182 22337
rect 17136 22265 17182 22303
rect 17136 22231 17142 22265
rect 17176 22231 17182 22265
rect 17136 22193 17182 22231
rect 17080 22159 17092 22170
rect 17022 22130 17092 22159
rect 17022 22078 17029 22130
rect 17081 22078 17092 22130
rect 17022 22040 17092 22078
rect 17136 22159 17142 22193
rect 17176 22159 17182 22193
rect 17232 23887 17238 23921
rect 17272 23887 17278 23921
rect 17313 24001 17383 24041
rect 17313 23949 17320 24001
rect 17372 23949 17383 24001
rect 17313 23921 17383 23949
rect 17313 23911 17334 23921
rect 17232 23849 17278 23887
rect 17232 23815 17238 23849
rect 17272 23815 17278 23849
rect 17232 23777 17278 23815
rect 17232 23743 17238 23777
rect 17272 23743 17278 23777
rect 17232 23705 17278 23743
rect 17232 23671 17238 23705
rect 17272 23671 17278 23705
rect 17232 23633 17278 23671
rect 17232 23599 17238 23633
rect 17272 23599 17278 23633
rect 17232 23561 17278 23599
rect 17232 23527 17238 23561
rect 17272 23527 17278 23561
rect 17232 23489 17278 23527
rect 17232 23455 17238 23489
rect 17272 23455 17278 23489
rect 17232 23417 17278 23455
rect 17232 23383 17238 23417
rect 17272 23383 17278 23417
rect 17232 23345 17278 23383
rect 17232 23311 17238 23345
rect 17272 23311 17278 23345
rect 17232 23273 17278 23311
rect 17232 23239 17238 23273
rect 17272 23239 17278 23273
rect 17232 23201 17278 23239
rect 17232 23167 17238 23201
rect 17272 23167 17278 23201
rect 17232 23129 17278 23167
rect 17232 23095 17238 23129
rect 17272 23095 17278 23129
rect 17232 23057 17278 23095
rect 17232 23023 17238 23057
rect 17272 23023 17278 23057
rect 17232 22985 17278 23023
rect 17232 22951 17238 22985
rect 17272 22951 17278 22985
rect 17232 22913 17278 22951
rect 17232 22879 17238 22913
rect 17272 22879 17278 22913
rect 17232 22841 17278 22879
rect 17232 22807 17238 22841
rect 17272 22807 17278 22841
rect 17232 22769 17278 22807
rect 17232 22735 17238 22769
rect 17272 22735 17278 22769
rect 17232 22697 17278 22735
rect 17232 22663 17238 22697
rect 17272 22663 17278 22697
rect 17232 22625 17278 22663
rect 17232 22591 17238 22625
rect 17272 22591 17278 22625
rect 17232 22553 17278 22591
rect 17232 22519 17238 22553
rect 17272 22519 17278 22553
rect 17232 22481 17278 22519
rect 17232 22447 17238 22481
rect 17272 22447 17278 22481
rect 17232 22409 17278 22447
rect 17232 22375 17238 22409
rect 17272 22375 17278 22409
rect 17232 22337 17278 22375
rect 17232 22303 17238 22337
rect 17272 22303 17278 22337
rect 17232 22265 17278 22303
rect 17232 22231 17238 22265
rect 17272 22231 17278 22265
rect 17232 22193 17278 22231
rect 17232 22173 17238 22193
rect 17136 22121 17182 22159
rect 17136 22087 17142 22121
rect 17176 22087 17182 22121
rect 17136 22040 17182 22087
rect 17213 22159 17238 22173
rect 17272 22173 17278 22193
rect 17328 23887 17334 23911
rect 17368 23911 17383 23921
rect 17424 23993 17470 24040
rect 17424 23959 17430 23993
rect 17464 23959 17470 23993
rect 17424 23921 17470 23959
rect 17368 23887 17374 23911
rect 17328 23849 17374 23887
rect 17328 23815 17334 23849
rect 17368 23815 17374 23849
rect 17328 23777 17374 23815
rect 17328 23743 17334 23777
rect 17368 23743 17374 23777
rect 17328 23705 17374 23743
rect 17328 23671 17334 23705
rect 17368 23671 17374 23705
rect 17328 23633 17374 23671
rect 17328 23599 17334 23633
rect 17368 23599 17374 23633
rect 17328 23561 17374 23599
rect 17328 23527 17334 23561
rect 17368 23527 17374 23561
rect 17328 23489 17374 23527
rect 17328 23455 17334 23489
rect 17368 23455 17374 23489
rect 17328 23417 17374 23455
rect 17328 23383 17334 23417
rect 17368 23383 17374 23417
rect 17328 23345 17374 23383
rect 17328 23311 17334 23345
rect 17368 23311 17374 23345
rect 17328 23273 17374 23311
rect 17328 23239 17334 23273
rect 17368 23239 17374 23273
rect 17328 23201 17374 23239
rect 17328 23167 17334 23201
rect 17368 23167 17374 23201
rect 17328 23129 17374 23167
rect 17328 23095 17334 23129
rect 17368 23095 17374 23129
rect 17328 23057 17374 23095
rect 17328 23023 17334 23057
rect 17368 23023 17374 23057
rect 17328 22985 17374 23023
rect 17328 22951 17334 22985
rect 17368 22951 17374 22985
rect 17328 22913 17374 22951
rect 17328 22879 17334 22913
rect 17368 22879 17374 22913
rect 17328 22841 17374 22879
rect 17328 22807 17334 22841
rect 17368 22807 17374 22841
rect 17328 22769 17374 22807
rect 17328 22735 17334 22769
rect 17368 22735 17374 22769
rect 17328 22697 17374 22735
rect 17328 22663 17334 22697
rect 17368 22663 17374 22697
rect 17328 22625 17374 22663
rect 17328 22591 17334 22625
rect 17368 22591 17374 22625
rect 17328 22553 17374 22591
rect 17328 22519 17334 22553
rect 17368 22519 17374 22553
rect 17328 22481 17374 22519
rect 17328 22447 17334 22481
rect 17368 22447 17374 22481
rect 17328 22409 17374 22447
rect 17328 22375 17334 22409
rect 17368 22375 17374 22409
rect 17328 22337 17374 22375
rect 17328 22303 17334 22337
rect 17368 22303 17374 22337
rect 17328 22265 17374 22303
rect 17328 22231 17334 22265
rect 17368 22231 17374 22265
rect 17328 22193 17374 22231
rect 17272 22159 17283 22173
rect 17213 22133 17283 22159
rect 17213 22081 17220 22133
rect 17272 22081 17283 22133
rect 17213 22043 17283 22081
rect 17328 22159 17334 22193
rect 17368 22159 17374 22193
rect 17424 23887 17430 23921
rect 17464 23887 17470 23921
rect 17513 24001 17583 24041
rect 17513 23949 17520 24001
rect 17572 23949 17583 24001
rect 17513 23921 17583 23949
rect 17513 23911 17526 23921
rect 17424 23849 17470 23887
rect 17424 23815 17430 23849
rect 17464 23815 17470 23849
rect 17424 23777 17470 23815
rect 17424 23743 17430 23777
rect 17464 23743 17470 23777
rect 17424 23705 17470 23743
rect 17424 23671 17430 23705
rect 17464 23671 17470 23705
rect 17424 23633 17470 23671
rect 17424 23599 17430 23633
rect 17464 23599 17470 23633
rect 17424 23561 17470 23599
rect 17424 23527 17430 23561
rect 17464 23527 17470 23561
rect 17424 23489 17470 23527
rect 17424 23455 17430 23489
rect 17464 23455 17470 23489
rect 17424 23417 17470 23455
rect 17424 23383 17430 23417
rect 17464 23383 17470 23417
rect 17424 23345 17470 23383
rect 17424 23311 17430 23345
rect 17464 23311 17470 23345
rect 17424 23273 17470 23311
rect 17424 23239 17430 23273
rect 17464 23239 17470 23273
rect 17424 23201 17470 23239
rect 17424 23167 17430 23201
rect 17464 23167 17470 23201
rect 17424 23129 17470 23167
rect 17424 23095 17430 23129
rect 17464 23095 17470 23129
rect 17424 23057 17470 23095
rect 17424 23023 17430 23057
rect 17464 23023 17470 23057
rect 17424 22985 17470 23023
rect 17424 22951 17430 22985
rect 17464 22951 17470 22985
rect 17424 22913 17470 22951
rect 17424 22879 17430 22913
rect 17464 22879 17470 22913
rect 17424 22841 17470 22879
rect 17424 22807 17430 22841
rect 17464 22807 17470 22841
rect 17424 22769 17470 22807
rect 17424 22735 17430 22769
rect 17464 22735 17470 22769
rect 17424 22697 17470 22735
rect 17424 22663 17430 22697
rect 17464 22663 17470 22697
rect 17424 22625 17470 22663
rect 17424 22591 17430 22625
rect 17464 22591 17470 22625
rect 17424 22553 17470 22591
rect 17424 22519 17430 22553
rect 17464 22519 17470 22553
rect 17424 22481 17470 22519
rect 17424 22447 17430 22481
rect 17464 22447 17470 22481
rect 17424 22409 17470 22447
rect 17424 22375 17430 22409
rect 17464 22375 17470 22409
rect 17424 22337 17470 22375
rect 17424 22303 17430 22337
rect 17464 22303 17470 22337
rect 17424 22265 17470 22303
rect 17424 22231 17430 22265
rect 17464 22231 17470 22265
rect 17424 22193 17470 22231
rect 17424 22171 17430 22193
rect 17328 22121 17374 22159
rect 17328 22087 17334 22121
rect 17368 22087 17374 22121
rect 17232 22040 17278 22043
rect 17328 22040 17374 22087
rect 17412 22159 17430 22171
rect 17464 22171 17470 22193
rect 17520 23887 17526 23911
rect 17560 23911 17583 23921
rect 17616 23993 17662 24040
rect 17616 23959 17622 23993
rect 17656 23959 17662 23993
rect 17616 23921 17662 23959
rect 17560 23887 17566 23911
rect 17520 23849 17566 23887
rect 17520 23815 17526 23849
rect 17560 23815 17566 23849
rect 17520 23777 17566 23815
rect 17520 23743 17526 23777
rect 17560 23743 17566 23777
rect 17520 23705 17566 23743
rect 17520 23671 17526 23705
rect 17560 23671 17566 23705
rect 17520 23633 17566 23671
rect 17520 23599 17526 23633
rect 17560 23599 17566 23633
rect 17520 23561 17566 23599
rect 17520 23527 17526 23561
rect 17560 23527 17566 23561
rect 17520 23489 17566 23527
rect 17520 23455 17526 23489
rect 17560 23455 17566 23489
rect 17520 23417 17566 23455
rect 17520 23383 17526 23417
rect 17560 23383 17566 23417
rect 17520 23345 17566 23383
rect 17520 23311 17526 23345
rect 17560 23311 17566 23345
rect 17520 23273 17566 23311
rect 17520 23239 17526 23273
rect 17560 23239 17566 23273
rect 17520 23201 17566 23239
rect 17520 23167 17526 23201
rect 17560 23167 17566 23201
rect 17520 23129 17566 23167
rect 17520 23095 17526 23129
rect 17560 23095 17566 23129
rect 17520 23057 17566 23095
rect 17520 23023 17526 23057
rect 17560 23023 17566 23057
rect 17520 22985 17566 23023
rect 17520 22951 17526 22985
rect 17560 22951 17566 22985
rect 17520 22913 17566 22951
rect 17520 22879 17526 22913
rect 17560 22879 17566 22913
rect 17520 22841 17566 22879
rect 17520 22807 17526 22841
rect 17560 22807 17566 22841
rect 17520 22769 17566 22807
rect 17520 22735 17526 22769
rect 17560 22735 17566 22769
rect 17520 22697 17566 22735
rect 17520 22663 17526 22697
rect 17560 22663 17566 22697
rect 17520 22625 17566 22663
rect 17520 22591 17526 22625
rect 17560 22591 17566 22625
rect 17520 22553 17566 22591
rect 17520 22519 17526 22553
rect 17560 22519 17566 22553
rect 17520 22481 17566 22519
rect 17520 22447 17526 22481
rect 17560 22447 17566 22481
rect 17520 22409 17566 22447
rect 17520 22375 17526 22409
rect 17560 22375 17566 22409
rect 17520 22337 17566 22375
rect 17520 22303 17526 22337
rect 17560 22303 17566 22337
rect 17520 22265 17566 22303
rect 17520 22231 17526 22265
rect 17560 22231 17566 22265
rect 17520 22193 17566 22231
rect 17464 22159 17482 22171
rect 17412 22131 17482 22159
rect 17412 22079 17419 22131
rect 17471 22079 17482 22131
rect 17412 22041 17482 22079
rect 17520 22159 17526 22193
rect 17560 22159 17566 22193
rect 17616 23887 17622 23921
rect 17656 23887 17662 23921
rect 17616 23849 17662 23887
rect 17616 23815 17622 23849
rect 17656 23815 17662 23849
rect 17616 23777 17662 23815
rect 17616 23743 17622 23777
rect 17656 23743 17662 23777
rect 17616 23705 17662 23743
rect 17616 23671 17622 23705
rect 17656 23671 17662 23705
rect 17616 23633 17662 23671
rect 17616 23599 17622 23633
rect 17656 23599 17662 23633
rect 17616 23561 17662 23599
rect 17616 23527 17622 23561
rect 17656 23527 17662 23561
rect 17616 23489 17662 23527
rect 17616 23455 17622 23489
rect 17656 23455 17662 23489
rect 17616 23417 17662 23455
rect 17616 23383 17622 23417
rect 17656 23383 17662 23417
rect 17616 23345 17662 23383
rect 17616 23311 17622 23345
rect 17656 23311 17662 23345
rect 17616 23273 17662 23311
rect 17616 23239 17622 23273
rect 17656 23239 17662 23273
rect 17616 23201 17662 23239
rect 17616 23167 17622 23201
rect 17656 23167 17662 23201
rect 17616 23129 17662 23167
rect 17616 23095 17622 23129
rect 17656 23095 17662 23129
rect 17616 23057 17662 23095
rect 17616 23023 17622 23057
rect 17656 23023 17662 23057
rect 17616 22985 17662 23023
rect 17616 22951 17622 22985
rect 17656 22951 17662 22985
rect 17616 22913 17662 22951
rect 17616 22879 17622 22913
rect 17656 22879 17662 22913
rect 17616 22841 17662 22879
rect 17616 22807 17622 22841
rect 17656 22807 17662 22841
rect 17616 22769 17662 22807
rect 17616 22735 17622 22769
rect 17656 22735 17662 22769
rect 17616 22697 17662 22735
rect 17616 22663 17622 22697
rect 17656 22663 17662 22697
rect 17616 22625 17662 22663
rect 17616 22591 17622 22625
rect 17656 22591 17662 22625
rect 17616 22553 17662 22591
rect 17616 22519 17622 22553
rect 17656 22519 17662 22553
rect 17616 22481 17662 22519
rect 17616 22447 17622 22481
rect 17656 22447 17662 22481
rect 17616 22409 17662 22447
rect 17616 22375 17622 22409
rect 17656 22375 17662 22409
rect 17616 22337 17662 22375
rect 17616 22303 17622 22337
rect 17656 22303 17662 22337
rect 17616 22265 17662 22303
rect 17616 22231 17622 22265
rect 17656 22231 17662 22265
rect 17616 22193 17662 22231
rect 17616 22172 17622 22193
rect 17520 22121 17566 22159
rect 17520 22087 17526 22121
rect 17560 22087 17566 22121
rect 17424 22040 17470 22041
rect 17520 22040 17566 22087
rect 17603 22159 17622 22172
rect 17656 22172 17662 22193
rect 17656 22159 17673 22172
rect 17603 22132 17673 22159
rect 17603 22080 17610 22132
rect 17662 22080 17673 22132
rect 17603 22042 17673 22080
rect 17616 22040 17662 22042
rect 16112 21990 16158 22028
rect 16112 21956 16118 21990
rect 16152 21956 16158 21990
rect 16112 21918 16158 21956
rect 16690 22002 17530 22010
rect 16690 21968 16710 22002
rect 16744 21968 16902 22002
rect 16936 21968 17094 22002
rect 17128 21968 17286 22002
rect 17320 21968 17478 22002
rect 17512 21968 17530 22002
rect 16690 21940 17530 21968
rect 16112 21884 16118 21918
rect 16152 21884 16158 21918
rect 16112 21846 16158 21884
rect 16112 21812 16118 21846
rect 16152 21812 16158 21846
rect 16112 21774 16158 21812
rect 16112 21740 16118 21774
rect 16152 21740 16158 21774
rect 16112 21702 16158 21740
rect 16112 21668 16118 21702
rect 16152 21668 16158 21702
rect 16112 21630 16158 21668
rect 16112 21596 16118 21630
rect 16152 21596 16158 21630
rect 16112 21558 16158 21596
rect 16112 21524 16118 21558
rect 16152 21524 16158 21558
rect 16112 21486 16158 21524
rect 16112 21452 16118 21486
rect 16152 21452 16158 21486
rect 16112 21414 16158 21452
rect 16112 21380 16118 21414
rect 16152 21380 16158 21414
rect 16112 21342 16158 21380
rect 17350 21718 17530 21770
rect 17350 21612 17387 21718
rect 17493 21612 17530 21718
rect 17350 21370 17530 21612
rect 17390 21350 17480 21370
rect 16056 21308 16071 21311
rect 16001 21277 16071 21308
rect 16001 21225 16010 21277
rect 16062 21225 16071 21277
rect 16001 21191 16071 21225
rect 16112 21308 16118 21342
rect 16152 21308 16158 21342
rect 16112 21270 16158 21308
rect 16112 21236 16118 21270
rect 16152 21236 16158 21270
rect 16016 21189 16062 21191
rect 16112 21189 16158 21236
rect 16780 21330 17130 21350
rect 16780 21296 16804 21330
rect 16838 21313 17130 21330
rect 16838 21296 16877 21313
rect 16780 21258 16877 21296
rect 16780 21224 16804 21258
rect 16838 21224 16877 21258
rect 14732 21150 14778 21151
rect 15290 21145 15324 21179
rect 15358 21150 15390 21179
rect 16780 21186 16877 21224
rect 16780 21152 16804 21186
rect 16838 21152 16877 21186
rect 15358 21145 16120 21150
rect 15290 21142 16120 21145
rect 13710 21112 14650 21120
rect 13710 21078 14018 21112
rect 14052 21078 14210 21112
rect 14244 21078 14402 21112
rect 14436 21078 14594 21112
rect 14628 21078 14650 21112
rect 15290 21108 15878 21142
rect 15912 21108 16070 21142
rect 16104 21108 16120 21142
rect 15290 21080 16120 21108
rect 16780 21114 16877 21152
rect 16780 21080 16804 21114
rect 16838 21080 16877 21114
rect 13000 16224 13120 21070
rect 13710 21040 14650 21078
rect 16780 21042 16877 21080
rect 16780 21008 16804 21042
rect 16838 21008 16877 21042
rect 16780 20970 16877 21008
rect 16780 20936 16804 20970
rect 16838 20941 16877 20970
rect 16993 20941 17130 21313
rect 17390 21316 17414 21350
rect 17448 21316 17480 21350
rect 17390 21278 17480 21316
rect 17390 21244 17414 21278
rect 17448 21244 17480 21278
rect 17390 21206 17480 21244
rect 17390 21172 17414 21206
rect 17448 21172 17480 21206
rect 17390 21134 17480 21172
rect 17390 21100 17414 21134
rect 17448 21100 17480 21134
rect 17390 21070 17480 21100
rect 17406 21062 17456 21070
rect 17406 21028 17414 21062
rect 17448 21028 17456 21062
rect 17406 20990 17456 21028
rect 17406 20956 17414 20990
rect 17448 20956 17456 20990
rect 17406 20943 17456 20956
rect 16838 20936 17130 20941
rect 16780 20910 17130 20936
rect 14880 20546 15490 20570
rect 14880 20494 14940 20546
rect 14992 20518 15004 20546
rect 15056 20494 15068 20546
rect 15120 20494 15132 20546
rect 15184 20518 15196 20546
rect 15248 20494 15260 20546
rect 15312 20494 15324 20546
rect 15376 20518 15388 20546
rect 15440 20494 15490 20546
rect 14880 20484 14974 20494
rect 15008 20484 15166 20494
rect 15200 20484 15358 20494
rect 15392 20484 15490 20494
rect 14880 20480 15490 20484
rect 14962 20478 15020 20480
rect 15154 20478 15212 20480
rect 15346 20478 15404 20480
rect 14824 20432 14870 20446
rect 14920 20440 14966 20446
rect 14824 20398 14830 20432
rect 14864 20398 14870 20432
rect 14824 20360 14870 20398
rect 14824 20326 14830 20360
rect 14864 20326 14870 20360
rect 14824 20288 14870 20326
rect 14900 20432 14980 20440
rect 14900 20401 14926 20432
rect 14960 20401 14980 20432
rect 14900 20349 14914 20401
rect 14966 20349 14980 20401
rect 14900 20326 14926 20349
rect 14960 20326 14980 20349
rect 14900 20310 14980 20326
rect 15016 20432 15062 20446
rect 15112 20440 15158 20446
rect 15016 20398 15022 20432
rect 15056 20398 15062 20432
rect 15016 20360 15062 20398
rect 15016 20326 15022 20360
rect 15056 20326 15062 20360
rect 14824 20254 14830 20288
rect 14864 20254 14870 20288
rect 14824 20216 14870 20254
rect 14824 20182 14830 20216
rect 14864 20182 14870 20216
rect 14824 20144 14870 20182
rect 14824 20110 14830 20144
rect 14864 20110 14870 20144
rect 14824 20072 14870 20110
rect 14824 20038 14830 20072
rect 14864 20038 14870 20072
rect 14824 20000 14870 20038
rect 14824 19966 14830 20000
rect 14864 19966 14870 20000
rect 14824 19928 14870 19966
rect 14824 19894 14830 19928
rect 14864 19894 14870 19928
rect 14824 19856 14870 19894
rect 14824 19822 14830 19856
rect 14864 19822 14870 19856
rect 14824 19784 14870 19822
rect 14824 19750 14830 19784
rect 14864 19750 14870 19784
rect 13306 19720 13486 19734
rect 14136 19720 14316 19734
rect 13306 19714 13739 19720
rect 13306 19608 13331 19714
rect 13725 19608 13739 19714
rect 13306 19602 13739 19608
rect 13887 19714 14316 19720
rect 13887 19608 13900 19714
rect 14294 19608 14316 19714
rect 13887 19602 14316 19608
rect 13306 19334 13486 19602
rect 14136 19334 14316 19602
rect 13306 19328 13739 19334
rect 13306 19222 13331 19328
rect 13725 19222 13739 19328
rect 13306 19216 13739 19222
rect 13887 19328 14316 19334
rect 13887 19222 13900 19328
rect 14294 19222 14316 19328
rect 14824 19712 14870 19750
rect 14824 19678 14830 19712
rect 14864 19678 14870 19712
rect 14824 19640 14870 19678
rect 14824 19606 14830 19640
rect 14864 19606 14870 19640
rect 14824 19568 14870 19606
rect 14824 19534 14830 19568
rect 14864 19534 14870 19568
rect 14824 19496 14870 19534
rect 14824 19462 14830 19496
rect 14864 19462 14870 19496
rect 14824 19424 14870 19462
rect 14824 19390 14830 19424
rect 14864 19390 14870 19424
rect 14824 19352 14870 19390
rect 14824 19318 14830 19352
rect 14864 19318 14870 19352
rect 14824 19300 14870 19318
rect 14920 20288 14966 20310
rect 14920 20254 14926 20288
rect 14960 20254 14966 20288
rect 14920 20216 14966 20254
rect 14920 20182 14926 20216
rect 14960 20182 14966 20216
rect 14920 20144 14966 20182
rect 14920 20110 14926 20144
rect 14960 20110 14966 20144
rect 14920 20072 14966 20110
rect 14920 20038 14926 20072
rect 14960 20038 14966 20072
rect 14920 20000 14966 20038
rect 14920 19966 14926 20000
rect 14960 19966 14966 20000
rect 14920 19928 14966 19966
rect 14920 19894 14926 19928
rect 14960 19894 14966 19928
rect 14920 19856 14966 19894
rect 14920 19822 14926 19856
rect 14960 19822 14966 19856
rect 14920 19784 14966 19822
rect 14920 19750 14926 19784
rect 14960 19750 14966 19784
rect 14920 19712 14966 19750
rect 14920 19678 14926 19712
rect 14960 19678 14966 19712
rect 14920 19640 14966 19678
rect 14920 19606 14926 19640
rect 14960 19606 14966 19640
rect 14920 19568 14966 19606
rect 14920 19534 14926 19568
rect 14960 19534 14966 19568
rect 14920 19496 14966 19534
rect 14920 19462 14926 19496
rect 14960 19462 14966 19496
rect 14920 19424 14966 19462
rect 14920 19390 14926 19424
rect 14960 19390 14966 19424
rect 14920 19352 14966 19390
rect 14920 19318 14926 19352
rect 14960 19318 14966 19352
rect 13887 19216 14316 19222
rect 13306 18948 13486 19216
rect 14136 18948 14316 19216
rect 14810 19280 14890 19300
rect 14810 19261 14830 19280
rect 14864 19261 14890 19280
rect 14810 19209 14824 19261
rect 14876 19209 14890 19261
rect 14810 19208 14890 19209
rect 14810 19174 14830 19208
rect 14864 19174 14890 19208
rect 14810 19170 14890 19174
rect 14920 19280 14966 19318
rect 15016 20288 15062 20326
rect 15090 20432 15170 20440
rect 15090 20401 15118 20432
rect 15152 20401 15170 20432
rect 15090 20349 15104 20401
rect 15156 20349 15170 20401
rect 15090 20326 15118 20349
rect 15152 20326 15170 20349
rect 15090 20310 15170 20326
rect 15208 20432 15254 20446
rect 15304 20440 15350 20446
rect 15208 20398 15214 20432
rect 15248 20398 15254 20432
rect 15208 20360 15254 20398
rect 15208 20326 15214 20360
rect 15248 20326 15254 20360
rect 15016 20254 15022 20288
rect 15056 20254 15062 20288
rect 15016 20216 15062 20254
rect 15016 20182 15022 20216
rect 15056 20182 15062 20216
rect 15016 20144 15062 20182
rect 15016 20110 15022 20144
rect 15056 20110 15062 20144
rect 15016 20072 15062 20110
rect 15016 20038 15022 20072
rect 15056 20038 15062 20072
rect 15016 20000 15062 20038
rect 15016 19966 15022 20000
rect 15056 19966 15062 20000
rect 15016 19928 15062 19966
rect 15016 19894 15022 19928
rect 15056 19894 15062 19928
rect 15016 19856 15062 19894
rect 15016 19822 15022 19856
rect 15056 19822 15062 19856
rect 15016 19784 15062 19822
rect 15016 19750 15022 19784
rect 15056 19750 15062 19784
rect 15016 19712 15062 19750
rect 15016 19678 15022 19712
rect 15056 19678 15062 19712
rect 15016 19640 15062 19678
rect 15016 19606 15022 19640
rect 15056 19606 15062 19640
rect 15016 19568 15062 19606
rect 15016 19534 15022 19568
rect 15056 19534 15062 19568
rect 15016 19496 15062 19534
rect 15016 19462 15022 19496
rect 15056 19462 15062 19496
rect 15016 19424 15062 19462
rect 15016 19390 15022 19424
rect 15056 19390 15062 19424
rect 15016 19352 15062 19390
rect 15016 19318 15022 19352
rect 15056 19318 15062 19352
rect 15016 19300 15062 19318
rect 15112 20288 15158 20310
rect 15112 20254 15118 20288
rect 15152 20254 15158 20288
rect 15112 20216 15158 20254
rect 15112 20182 15118 20216
rect 15152 20182 15158 20216
rect 15112 20144 15158 20182
rect 15112 20110 15118 20144
rect 15152 20110 15158 20144
rect 15112 20072 15158 20110
rect 15112 20038 15118 20072
rect 15152 20038 15158 20072
rect 15112 20000 15158 20038
rect 15112 19966 15118 20000
rect 15152 19966 15158 20000
rect 15112 19928 15158 19966
rect 15112 19894 15118 19928
rect 15152 19894 15158 19928
rect 15112 19856 15158 19894
rect 15112 19822 15118 19856
rect 15152 19822 15158 19856
rect 15112 19784 15158 19822
rect 15112 19750 15118 19784
rect 15152 19750 15158 19784
rect 15112 19712 15158 19750
rect 15112 19678 15118 19712
rect 15152 19678 15158 19712
rect 15112 19640 15158 19678
rect 15112 19606 15118 19640
rect 15152 19606 15158 19640
rect 15112 19568 15158 19606
rect 15112 19534 15118 19568
rect 15152 19534 15158 19568
rect 15112 19496 15158 19534
rect 15112 19462 15118 19496
rect 15152 19462 15158 19496
rect 15112 19424 15158 19462
rect 15112 19390 15118 19424
rect 15152 19390 15158 19424
rect 15112 19352 15158 19390
rect 15112 19318 15118 19352
rect 15152 19318 15158 19352
rect 14920 19246 14926 19280
rect 14960 19246 14966 19280
rect 14920 19208 14966 19246
rect 14920 19174 14926 19208
rect 14960 19174 14966 19208
rect 14824 19160 14870 19170
rect 14920 19160 14966 19174
rect 15000 19280 15080 19300
rect 15000 19261 15022 19280
rect 15056 19261 15080 19280
rect 15000 19209 15014 19261
rect 15066 19209 15080 19261
rect 15000 19208 15080 19209
rect 15000 19174 15022 19208
rect 15056 19174 15080 19208
rect 15000 19170 15080 19174
rect 15112 19280 15158 19318
rect 15208 20288 15254 20326
rect 15290 20432 15370 20440
rect 15290 20401 15310 20432
rect 15344 20401 15370 20432
rect 15290 20349 15304 20401
rect 15356 20349 15370 20401
rect 15290 20326 15310 20349
rect 15344 20326 15370 20349
rect 15290 20310 15370 20326
rect 15400 20432 15446 20446
rect 15496 20440 15542 20446
rect 15400 20398 15406 20432
rect 15440 20398 15446 20432
rect 15400 20360 15446 20398
rect 15400 20326 15406 20360
rect 15440 20326 15446 20360
rect 15208 20254 15214 20288
rect 15248 20254 15254 20288
rect 15208 20216 15254 20254
rect 15208 20182 15214 20216
rect 15248 20182 15254 20216
rect 15208 20144 15254 20182
rect 15208 20110 15214 20144
rect 15248 20110 15254 20144
rect 15208 20072 15254 20110
rect 15208 20038 15214 20072
rect 15248 20038 15254 20072
rect 15208 20000 15254 20038
rect 15208 19966 15214 20000
rect 15248 19966 15254 20000
rect 15208 19928 15254 19966
rect 15208 19894 15214 19928
rect 15248 19894 15254 19928
rect 15208 19856 15254 19894
rect 15208 19822 15214 19856
rect 15248 19822 15254 19856
rect 15208 19784 15254 19822
rect 15208 19750 15214 19784
rect 15248 19750 15254 19784
rect 15208 19712 15254 19750
rect 15208 19678 15214 19712
rect 15248 19678 15254 19712
rect 15208 19640 15254 19678
rect 15208 19606 15214 19640
rect 15248 19606 15254 19640
rect 15208 19568 15254 19606
rect 15208 19534 15214 19568
rect 15248 19534 15254 19568
rect 15208 19496 15254 19534
rect 15208 19462 15214 19496
rect 15248 19462 15254 19496
rect 15208 19424 15254 19462
rect 15208 19390 15214 19424
rect 15248 19390 15254 19424
rect 15208 19352 15254 19390
rect 15208 19318 15214 19352
rect 15248 19318 15254 19352
rect 15208 19300 15254 19318
rect 15304 20288 15350 20310
rect 15304 20254 15310 20288
rect 15344 20254 15350 20288
rect 15304 20216 15350 20254
rect 15304 20182 15310 20216
rect 15344 20182 15350 20216
rect 15304 20144 15350 20182
rect 15304 20110 15310 20144
rect 15344 20110 15350 20144
rect 15304 20072 15350 20110
rect 15304 20038 15310 20072
rect 15344 20038 15350 20072
rect 15304 20000 15350 20038
rect 15304 19966 15310 20000
rect 15344 19966 15350 20000
rect 15304 19928 15350 19966
rect 15304 19894 15310 19928
rect 15344 19894 15350 19928
rect 15304 19856 15350 19894
rect 15304 19822 15310 19856
rect 15344 19822 15350 19856
rect 15304 19784 15350 19822
rect 15304 19750 15310 19784
rect 15344 19750 15350 19784
rect 15304 19712 15350 19750
rect 15304 19678 15310 19712
rect 15344 19678 15350 19712
rect 15304 19640 15350 19678
rect 15304 19606 15310 19640
rect 15344 19606 15350 19640
rect 15304 19568 15350 19606
rect 15304 19534 15310 19568
rect 15344 19534 15350 19568
rect 15304 19496 15350 19534
rect 15304 19462 15310 19496
rect 15344 19462 15350 19496
rect 15304 19424 15350 19462
rect 15304 19390 15310 19424
rect 15344 19390 15350 19424
rect 15304 19352 15350 19390
rect 15304 19318 15310 19352
rect 15344 19318 15350 19352
rect 15112 19246 15118 19280
rect 15152 19246 15158 19280
rect 15112 19208 15158 19246
rect 15112 19174 15118 19208
rect 15152 19174 15158 19208
rect 15016 19160 15062 19170
rect 15112 19160 15158 19174
rect 15190 19280 15270 19300
rect 15190 19261 15214 19280
rect 15248 19261 15270 19280
rect 15190 19209 15204 19261
rect 15256 19209 15270 19261
rect 15190 19208 15270 19209
rect 15190 19174 15214 19208
rect 15248 19174 15270 19208
rect 15190 19170 15270 19174
rect 15304 19280 15350 19318
rect 15400 20288 15446 20326
rect 15480 20432 15560 20440
rect 15480 20401 15502 20432
rect 15536 20401 15560 20432
rect 15480 20349 15494 20401
rect 15546 20349 15560 20401
rect 15480 20326 15502 20349
rect 15536 20326 15560 20349
rect 15480 20310 15560 20326
rect 15400 20254 15406 20288
rect 15440 20254 15446 20288
rect 15400 20216 15446 20254
rect 15400 20182 15406 20216
rect 15440 20182 15446 20216
rect 15400 20144 15446 20182
rect 15400 20110 15406 20144
rect 15440 20110 15446 20144
rect 15400 20072 15446 20110
rect 15400 20038 15406 20072
rect 15440 20038 15446 20072
rect 15400 20000 15446 20038
rect 15400 19966 15406 20000
rect 15440 19966 15446 20000
rect 15400 19928 15446 19966
rect 15400 19894 15406 19928
rect 15440 19894 15446 19928
rect 15400 19856 15446 19894
rect 15400 19822 15406 19856
rect 15440 19822 15446 19856
rect 15400 19784 15446 19822
rect 15400 19750 15406 19784
rect 15440 19750 15446 19784
rect 15400 19712 15446 19750
rect 15400 19678 15406 19712
rect 15440 19678 15446 19712
rect 15400 19640 15446 19678
rect 15400 19606 15406 19640
rect 15440 19606 15446 19640
rect 15400 19568 15446 19606
rect 15400 19534 15406 19568
rect 15440 19534 15446 19568
rect 15400 19496 15446 19534
rect 15400 19462 15406 19496
rect 15440 19462 15446 19496
rect 15400 19424 15446 19462
rect 15400 19390 15406 19424
rect 15440 19390 15446 19424
rect 15400 19352 15446 19390
rect 15400 19318 15406 19352
rect 15440 19318 15446 19352
rect 15400 19300 15446 19318
rect 15496 20288 15542 20310
rect 15496 20254 15502 20288
rect 15536 20254 15542 20288
rect 15496 20216 15542 20254
rect 15496 20182 15502 20216
rect 15536 20182 15542 20216
rect 15496 20144 15542 20182
rect 15496 20110 15502 20144
rect 15536 20110 15542 20144
rect 15496 20072 15542 20110
rect 15496 20038 15502 20072
rect 15536 20038 15542 20072
rect 15496 20000 15542 20038
rect 15496 19966 15502 20000
rect 15536 19966 15542 20000
rect 16120 20032 16180 20050
rect 16120 19998 16134 20032
rect 16168 19998 16180 20032
rect 16120 19990 16180 19998
rect 15496 19928 15542 19966
rect 15496 19894 15502 19928
rect 15536 19894 15542 19928
rect 15496 19856 15542 19894
rect 15496 19822 15502 19856
rect 15536 19822 15542 19856
rect 15496 19784 15542 19822
rect 15496 19750 15502 19784
rect 15536 19750 15542 19784
rect 15496 19712 15542 19750
rect 15496 19678 15502 19712
rect 15536 19678 15542 19712
rect 15496 19640 15542 19678
rect 15496 19606 15502 19640
rect 15536 19606 15542 19640
rect 15496 19568 15542 19606
rect 15496 19534 15502 19568
rect 15536 19534 15542 19568
rect 15496 19496 15542 19534
rect 15496 19462 15502 19496
rect 15536 19462 15542 19496
rect 15496 19424 15542 19462
rect 15496 19390 15502 19424
rect 15536 19390 15542 19424
rect 15496 19352 15542 19390
rect 15496 19318 15502 19352
rect 15536 19318 15542 19352
rect 15304 19246 15310 19280
rect 15344 19246 15350 19280
rect 15304 19208 15350 19246
rect 15304 19174 15310 19208
rect 15344 19174 15350 19208
rect 15208 19160 15254 19170
rect 15304 19160 15350 19174
rect 15380 19280 15460 19300
rect 15380 19261 15406 19280
rect 15440 19261 15460 19280
rect 15380 19209 15394 19261
rect 15446 19209 15460 19261
rect 15380 19208 15460 19209
rect 15380 19174 15406 19208
rect 15440 19174 15460 19208
rect 15380 19170 15460 19174
rect 15496 19280 15542 19318
rect 15984 19937 16030 19960
rect 15984 19903 15990 19937
rect 16024 19903 16030 19937
rect 15984 19865 16030 19903
rect 15984 19831 15990 19865
rect 16024 19831 16030 19865
rect 15984 19793 16030 19831
rect 16060 19937 16140 19960
rect 16060 19921 16086 19937
rect 16120 19921 16140 19937
rect 16060 19869 16074 19921
rect 16126 19869 16140 19921
rect 16060 19865 16140 19869
rect 16060 19831 16086 19865
rect 16120 19831 16140 19865
rect 16060 19830 16140 19831
rect 16176 19937 16222 19960
rect 16176 19903 16182 19937
rect 16216 19903 16222 19937
rect 16176 19865 16222 19903
rect 16176 19831 16182 19865
rect 16216 19831 16222 19865
rect 15984 19759 15990 19793
rect 16024 19759 16030 19793
rect 15984 19721 16030 19759
rect 15984 19687 15990 19721
rect 16024 19687 16030 19721
rect 15984 19649 16030 19687
rect 15984 19615 15990 19649
rect 16024 19615 16030 19649
rect 15984 19577 16030 19615
rect 15984 19543 15990 19577
rect 16024 19543 16030 19577
rect 15984 19505 16030 19543
rect 15984 19471 15990 19505
rect 16024 19471 16030 19505
rect 15984 19433 16030 19471
rect 15984 19399 15990 19433
rect 16024 19399 16030 19433
rect 15984 19361 16030 19399
rect 15984 19327 15990 19361
rect 16024 19327 16030 19361
rect 15984 19290 16030 19327
rect 16080 19793 16126 19830
rect 16080 19759 16086 19793
rect 16120 19759 16126 19793
rect 16080 19721 16126 19759
rect 16080 19687 16086 19721
rect 16120 19687 16126 19721
rect 16080 19649 16126 19687
rect 16080 19615 16086 19649
rect 16120 19615 16126 19649
rect 16080 19577 16126 19615
rect 16080 19543 16086 19577
rect 16120 19543 16126 19577
rect 16080 19505 16126 19543
rect 16080 19471 16086 19505
rect 16120 19471 16126 19505
rect 16080 19433 16126 19471
rect 16080 19399 16086 19433
rect 16120 19399 16126 19433
rect 16080 19361 16126 19399
rect 16080 19327 16086 19361
rect 16120 19327 16126 19361
rect 15496 19246 15502 19280
rect 15536 19246 15542 19280
rect 15496 19208 15542 19246
rect 15496 19174 15502 19208
rect 15536 19174 15542 19208
rect 15400 19160 15446 19170
rect 15496 19160 15542 19174
rect 15960 19289 16040 19290
rect 15960 19255 15990 19289
rect 16024 19255 16040 19289
rect 15960 19251 16040 19255
rect 15960 19199 15974 19251
rect 16026 19199 16040 19251
rect 15960 19183 15990 19199
rect 16024 19183 16040 19199
rect 15960 19160 16040 19183
rect 16080 19289 16126 19327
rect 16176 19793 16222 19831
rect 16250 19937 16330 19960
rect 16250 19921 16278 19937
rect 16312 19921 16330 19937
rect 16250 19869 16264 19921
rect 16316 19869 16330 19921
rect 16250 19865 16330 19869
rect 16250 19831 16278 19865
rect 16312 19831 16330 19865
rect 16250 19830 16330 19831
rect 16176 19759 16182 19793
rect 16216 19759 16222 19793
rect 16176 19721 16222 19759
rect 16176 19687 16182 19721
rect 16216 19687 16222 19721
rect 16176 19649 16222 19687
rect 16176 19615 16182 19649
rect 16216 19615 16222 19649
rect 16176 19577 16222 19615
rect 16176 19543 16182 19577
rect 16216 19543 16222 19577
rect 16176 19505 16222 19543
rect 16176 19471 16182 19505
rect 16216 19471 16222 19505
rect 16176 19433 16222 19471
rect 16176 19399 16182 19433
rect 16216 19399 16222 19433
rect 16176 19361 16222 19399
rect 16176 19327 16182 19361
rect 16216 19327 16222 19361
rect 16176 19290 16222 19327
rect 16272 19793 16318 19830
rect 16272 19759 16278 19793
rect 16312 19759 16318 19793
rect 16272 19721 16318 19759
rect 16272 19687 16278 19721
rect 16312 19687 16318 19721
rect 16272 19649 16318 19687
rect 16272 19615 16278 19649
rect 16312 19615 16318 19649
rect 16272 19577 16318 19615
rect 16272 19543 16278 19577
rect 16312 19543 16318 19577
rect 16272 19505 16318 19543
rect 16272 19471 16278 19505
rect 16312 19471 16318 19505
rect 16272 19433 16318 19471
rect 16272 19399 16278 19433
rect 16312 19399 16318 19433
rect 16272 19361 16318 19399
rect 16272 19327 16278 19361
rect 16312 19327 16318 19361
rect 16080 19255 16086 19289
rect 16120 19255 16126 19289
rect 16080 19217 16126 19255
rect 16080 19183 16086 19217
rect 16120 19183 16126 19217
rect 16080 19160 16126 19183
rect 16160 19289 16240 19290
rect 16160 19255 16182 19289
rect 16216 19255 16240 19289
rect 16160 19251 16240 19255
rect 16160 19199 16174 19251
rect 16226 19199 16240 19251
rect 16160 19183 16182 19199
rect 16216 19183 16240 19199
rect 16160 19160 16240 19183
rect 16272 19289 16318 19327
rect 16272 19255 16278 19289
rect 16312 19255 16318 19289
rect 16272 19217 16318 19255
rect 16272 19183 16278 19217
rect 16312 19183 16318 19217
rect 16272 19160 16318 19183
rect 16796 19299 16846 19313
rect 16796 19265 16804 19299
rect 16838 19265 16846 19299
rect 16796 19227 16846 19265
rect 16796 19193 16804 19227
rect 16838 19193 16846 19227
rect 16796 19155 16846 19193
rect 17020 19241 17230 19280
rect 17020 19189 17067 19241
rect 17119 19189 17131 19241
rect 17183 19189 17230 19241
rect 17020 19160 17230 19189
rect 14860 19122 15510 19130
rect 14860 19088 14878 19122
rect 14912 19088 15070 19122
rect 15104 19088 15262 19122
rect 15296 19088 15454 19122
rect 15488 19088 15510 19122
rect 14860 19060 15510 19088
rect 16020 19122 16610 19130
rect 16020 19088 16038 19122
rect 16072 19088 16230 19122
rect 16264 19101 16610 19122
rect 16264 19088 16524 19101
rect 16020 19070 16524 19088
rect 13306 18942 13739 18948
rect 13306 18836 13331 18942
rect 13725 18836 13739 18942
rect 13306 18830 13739 18836
rect 13887 18942 14316 18948
rect 13887 18836 13900 18942
rect 14294 18836 14316 18942
rect 15140 18980 15260 19060
rect 16490 19049 16524 19070
rect 16576 19049 16610 19101
rect 16490 19020 16610 19049
rect 16796 19121 16804 19155
rect 16838 19121 16846 19155
rect 16796 19083 16846 19121
rect 16796 19049 16804 19083
rect 16838 19049 16846 19083
rect 16796 19011 16846 19049
rect 16796 18980 16804 19011
rect 15140 18977 16804 18980
rect 16838 18980 16846 19011
rect 16838 18977 16860 18980
rect 15140 18939 16860 18977
rect 15140 18905 16804 18939
rect 16838 18905 16860 18939
rect 15140 18860 16860 18905
rect 13887 18830 14316 18836
rect 13306 18562 13486 18830
rect 14136 18562 14316 18830
rect 15038 18714 16326 18787
rect 15038 18584 15111 18714
rect 13306 18556 13739 18562
rect 13306 18450 13331 18556
rect 13725 18450 13739 18556
rect 13306 18444 13739 18450
rect 13887 18556 14316 18562
rect 13887 18450 13900 18556
rect 14294 18450 14316 18556
rect 15036 18566 15116 18584
rect 15036 18532 15060 18566
rect 15094 18532 15116 18566
rect 15036 18524 15116 18532
rect 15446 18566 15526 18584
rect 15446 18532 15470 18566
rect 15504 18532 15526 18566
rect 15446 18524 15526 18532
rect 16253 18535 16326 18714
rect 16253 18501 16272 18535
rect 16306 18501 16326 18535
rect 13887 18444 14316 18450
rect 13306 18176 13486 18444
rect 14136 18176 14316 18444
rect 15010 18451 15056 18494
rect 15010 18417 15016 18451
rect 15050 18417 15056 18451
rect 15010 18379 15056 18417
rect 15010 18345 15016 18379
rect 15050 18345 15056 18379
rect 15010 18307 15056 18345
rect 15010 18273 15016 18307
rect 15050 18273 15056 18307
rect 15010 18235 15056 18273
rect 15010 18209 15016 18235
rect 13306 18170 13739 18176
rect 13306 18064 13331 18170
rect 13725 18064 13739 18170
rect 13306 18058 13739 18064
rect 13887 18170 14316 18176
rect 13887 18064 13900 18170
rect 14294 18064 14316 18170
rect 13887 18058 14316 18064
rect 13306 17790 13486 18058
rect 14136 17790 14316 18058
rect 13306 17784 13739 17790
rect 13306 17678 13331 17784
rect 13725 17678 13739 17784
rect 13306 17672 13739 17678
rect 13887 17784 14316 17790
rect 13887 17678 13900 17784
rect 14294 17678 14316 17784
rect 13887 17672 14316 17678
rect 13306 17404 13486 17672
rect 14136 17404 14316 17672
rect 13306 17398 13739 17404
rect 13306 17292 13331 17398
rect 13725 17292 13739 17398
rect 13306 17286 13739 17292
rect 13887 17398 14316 17404
rect 13887 17292 13900 17398
rect 14294 17292 14316 17398
rect 13887 17286 14316 17292
rect 13306 17018 13486 17286
rect 14136 17018 14316 17286
rect 13306 17012 13739 17018
rect 13306 16906 13331 17012
rect 13725 16906 13739 17012
rect 13306 16900 13739 16906
rect 13887 17012 14316 17018
rect 13887 16906 13900 17012
rect 14294 16906 14316 17012
rect 13887 16900 14316 16906
rect 13306 16432 13486 16900
rect 14136 16692 14316 16900
rect 14136 16576 14163 16692
rect 14279 16576 14316 16692
rect 14136 16554 14316 16576
rect 14371 18201 15016 18209
rect 15050 18201 15056 18235
rect 14371 18163 15056 18201
rect 14371 18129 15016 18163
rect 15050 18129 15056 18163
rect 14371 18096 15056 18129
rect 13306 16326 13338 16432
rect 13444 16326 13486 16432
rect 13306 16304 13486 16326
rect 13516 16392 13612 16397
rect 14371 16392 14484 18096
rect 15010 18091 15056 18096
rect 15010 18057 15016 18091
rect 15050 18057 15056 18091
rect 15010 18019 15056 18057
rect 15010 17985 15016 18019
rect 15050 17985 15056 18019
rect 15010 17947 15056 17985
rect 15010 17913 15016 17947
rect 15050 17913 15056 17947
rect 15010 17875 15056 17913
rect 14641 17834 14755 17851
rect 14641 17800 14660 17834
rect 14694 17809 14755 17834
rect 14641 17762 14669 17800
rect 14641 17728 14660 17762
rect 14721 17757 14755 17809
rect 14694 17745 14755 17757
rect 14641 17693 14669 17728
rect 14721 17693 14755 17745
rect 14641 17690 14755 17693
rect 14641 17656 14660 17690
rect 14694 17681 14755 17690
rect 14641 17629 14669 17656
rect 14721 17629 14755 17681
rect 14641 17618 14755 17629
rect 14641 17594 14660 17618
rect 14652 17584 14660 17594
rect 14694 17594 14755 17618
rect 15010 17841 15016 17875
rect 15050 17841 15056 17875
rect 15010 17803 15056 17841
rect 15010 17769 15016 17803
rect 15050 17769 15056 17803
rect 15010 17731 15056 17769
rect 15010 17697 15016 17731
rect 15050 17697 15056 17731
rect 15010 17659 15056 17697
rect 15010 17625 15016 17659
rect 15050 17625 15056 17659
rect 14694 17584 14702 17594
rect 14652 17546 14702 17584
rect 14652 17512 14660 17546
rect 14694 17512 14702 17546
rect 14652 17474 14702 17512
rect 14652 17440 14660 17474
rect 14694 17440 14702 17474
rect 14652 17427 14702 17440
rect 15010 17587 15056 17625
rect 15010 17553 15016 17587
rect 15050 17553 15056 17587
rect 15010 17515 15056 17553
rect 15010 17481 15016 17515
rect 15050 17481 15056 17515
rect 15010 17443 15056 17481
rect 15010 17409 15016 17443
rect 15050 17409 15056 17443
rect 15010 17371 15056 17409
rect 15010 17337 15016 17371
rect 15050 17337 15056 17371
rect 14652 17303 14702 17317
rect 14652 17269 14660 17303
rect 14694 17269 14702 17303
rect 14652 17231 14702 17269
rect 14652 17197 14660 17231
rect 14694 17197 14702 17231
rect 14652 17159 14702 17197
rect 14652 17125 14660 17159
rect 14694 17125 14702 17159
rect 14652 17087 14702 17125
rect 14652 17053 14660 17087
rect 14694 17053 14702 17087
rect 14652 17015 14702 17053
rect 14652 17004 14660 17015
rect 13516 16362 14484 16392
rect 13516 16310 13534 16362
rect 13586 16310 14484 16362
rect 14596 16981 14660 17004
rect 14694 17004 14702 17015
rect 15010 17299 15056 17337
rect 15010 17265 15016 17299
rect 15050 17265 15056 17299
rect 15010 17227 15056 17265
rect 15010 17193 15016 17227
rect 15050 17193 15056 17227
rect 15010 17155 15056 17193
rect 15010 17121 15016 17155
rect 15050 17121 15056 17155
rect 15010 17083 15056 17121
rect 15010 17049 15016 17083
rect 15050 17049 15056 17083
rect 15010 17011 15056 17049
rect 14694 16981 14756 17004
rect 14596 16943 14756 16981
rect 14596 16909 14660 16943
rect 14694 16909 14756 16943
rect 15010 16977 15016 17011
rect 15050 16977 15056 17011
rect 15010 16934 15056 16977
rect 15098 18451 15144 18494
rect 15098 18417 15104 18451
rect 15138 18417 15144 18451
rect 15098 18379 15144 18417
rect 15098 18345 15104 18379
rect 15138 18345 15144 18379
rect 15098 18307 15144 18345
rect 15098 18273 15104 18307
rect 15138 18273 15144 18307
rect 15098 18235 15144 18273
rect 15098 18201 15104 18235
rect 15138 18201 15144 18235
rect 15098 18163 15144 18201
rect 15098 18129 15104 18163
rect 15138 18129 15144 18163
rect 15098 18091 15144 18129
rect 15098 18057 15104 18091
rect 15138 18057 15144 18091
rect 15098 18019 15144 18057
rect 15098 17985 15104 18019
rect 15138 17985 15144 18019
rect 15098 17947 15144 17985
rect 15098 17913 15104 17947
rect 15138 17913 15144 17947
rect 15098 17875 15144 17913
rect 15098 17841 15104 17875
rect 15138 17851 15144 17875
rect 15420 18451 15466 18494
rect 15420 18417 15426 18451
rect 15460 18417 15466 18451
rect 15420 18379 15466 18417
rect 15420 18345 15426 18379
rect 15460 18345 15466 18379
rect 15420 18307 15466 18345
rect 15420 18273 15426 18307
rect 15460 18273 15466 18307
rect 15420 18235 15466 18273
rect 15420 18201 15426 18235
rect 15460 18201 15466 18235
rect 15420 18163 15466 18201
rect 15420 18129 15426 18163
rect 15460 18129 15466 18163
rect 15420 18091 15466 18129
rect 15420 18057 15426 18091
rect 15460 18057 15466 18091
rect 15420 18019 15466 18057
rect 15420 17985 15426 18019
rect 15460 17985 15466 18019
rect 15420 17947 15466 17985
rect 15420 17913 15426 17947
rect 15460 17913 15466 17947
rect 15420 17875 15466 17913
rect 15138 17841 15187 17851
rect 15098 17810 15187 17841
rect 15098 17803 15119 17810
rect 15098 17769 15104 17803
rect 15098 17758 15119 17769
rect 15171 17758 15187 17810
rect 15098 17746 15187 17758
rect 15098 17731 15119 17746
rect 15098 17697 15104 17731
rect 15098 17694 15119 17697
rect 15171 17694 15187 17746
rect 15098 17682 15187 17694
rect 15098 17659 15119 17682
rect 15098 17625 15104 17659
rect 15171 17630 15187 17682
rect 15138 17625 15187 17630
rect 15098 17596 15187 17625
rect 15420 17841 15426 17875
rect 15460 17841 15466 17875
rect 15508 18451 15554 18494
rect 15508 18417 15514 18451
rect 15548 18417 15554 18451
rect 15508 18379 15554 18417
rect 16253 18463 16326 18501
rect 16253 18429 16272 18463
rect 16306 18429 16326 18463
rect 16253 18409 16326 18429
rect 15508 18345 15514 18379
rect 15548 18345 15554 18379
rect 15508 18307 15554 18345
rect 15508 18273 15514 18307
rect 15548 18273 15554 18307
rect 15508 18235 15554 18273
rect 15508 18201 15514 18235
rect 15548 18201 15554 18235
rect 16264 18391 16314 18409
rect 16264 18357 16272 18391
rect 16306 18357 16314 18391
rect 16264 18319 16314 18357
rect 16788 18350 16878 18352
rect 16264 18285 16272 18319
rect 16306 18285 16314 18319
rect 16264 18247 16314 18285
rect 15508 18163 15554 18201
rect 15508 18129 15514 18163
rect 15548 18129 15554 18163
rect 15508 18091 15554 18129
rect 15508 18057 15514 18091
rect 15548 18057 15554 18091
rect 15508 18019 15554 18057
rect 15508 17985 15514 18019
rect 15548 17985 15554 18019
rect 15508 17947 15554 17985
rect 15508 17913 15514 17947
rect 15548 17913 15554 17947
rect 15508 17875 15554 17913
rect 15508 17857 15514 17875
rect 15420 17803 15466 17841
rect 15420 17769 15426 17803
rect 15460 17769 15466 17803
rect 15420 17731 15466 17769
rect 15420 17697 15426 17731
rect 15460 17697 15466 17731
rect 15420 17659 15466 17697
rect 15420 17625 15426 17659
rect 15460 17625 15466 17659
rect 15098 17587 15144 17596
rect 15098 17553 15104 17587
rect 15138 17553 15144 17587
rect 15098 17515 15144 17553
rect 15098 17481 15104 17515
rect 15138 17481 15144 17515
rect 15098 17443 15144 17481
rect 15098 17409 15104 17443
rect 15138 17409 15144 17443
rect 15098 17371 15144 17409
rect 15098 17337 15104 17371
rect 15138 17337 15144 17371
rect 15098 17299 15144 17337
rect 15098 17265 15104 17299
rect 15138 17265 15144 17299
rect 15098 17227 15144 17265
rect 15098 17193 15104 17227
rect 15138 17193 15144 17227
rect 15098 17155 15144 17193
rect 15098 17121 15104 17155
rect 15138 17121 15144 17155
rect 15098 17083 15144 17121
rect 15098 17049 15104 17083
rect 15138 17049 15144 17083
rect 15098 17044 15144 17049
rect 15420 17587 15466 17625
rect 15506 17841 15514 17857
rect 15548 17857 15554 17875
rect 15787 17870 15974 18232
rect 16264 18213 16272 18247
rect 16306 18213 16314 18247
rect 16264 18175 16314 18213
rect 16264 18141 16272 18175
rect 16306 18141 16314 18175
rect 16264 18128 16314 18141
rect 16780 18330 16880 18350
rect 16780 18296 16816 18330
rect 16850 18296 16880 18330
rect 16780 18016 16880 18296
rect 16780 17964 16804 18016
rect 16856 17964 16880 18016
rect 16780 17930 16880 17964
rect 17330 18012 17530 18060
rect 15780 17857 16980 17870
rect 15548 17841 16980 17857
rect 15506 17834 16980 17841
rect 15506 17803 15880 17834
rect 15506 17769 15514 17803
rect 15548 17800 15880 17803
rect 15914 17800 16980 17834
rect 15548 17769 16980 17800
rect 15506 17762 16980 17769
rect 15506 17731 15880 17762
rect 15506 17697 15514 17731
rect 15548 17728 15880 17731
rect 15914 17728 16980 17762
rect 15548 17697 16980 17728
rect 17330 17768 17372 18012
rect 17488 17768 17530 18012
rect 17330 17741 17414 17768
rect 17448 17741 17530 17768
rect 17330 17720 17530 17741
rect 15506 17690 16980 17697
rect 15506 17659 15880 17690
rect 15506 17625 15514 17659
rect 15548 17656 15880 17659
rect 15914 17656 16980 17690
rect 15548 17625 16980 17656
rect 15506 17618 16980 17625
rect 15506 17601 15880 17618
rect 15420 17553 15426 17587
rect 15460 17553 15466 17587
rect 15420 17515 15466 17553
rect 15420 17481 15426 17515
rect 15460 17481 15466 17515
rect 15420 17443 15466 17481
rect 15420 17409 15426 17443
rect 15460 17409 15466 17443
rect 15420 17371 15466 17409
rect 15420 17337 15426 17371
rect 15460 17337 15466 17371
rect 15420 17299 15466 17337
rect 15420 17265 15426 17299
rect 15460 17265 15466 17299
rect 15420 17227 15466 17265
rect 15420 17193 15426 17227
rect 15460 17193 15466 17227
rect 15420 17155 15466 17193
rect 15420 17121 15426 17155
rect 15460 17121 15466 17155
rect 15420 17083 15466 17121
rect 15420 17049 15426 17083
rect 15460 17049 15466 17083
rect 15098 17011 15265 17044
rect 15098 16977 15104 17011
rect 15138 16977 15265 17011
rect 15098 16943 15265 16977
rect 15420 17011 15466 17049
rect 15420 16977 15426 17011
rect 15460 16977 15466 17011
rect 15098 16934 15144 16943
rect 15420 16934 15466 16977
rect 15508 17587 15554 17601
rect 15508 17553 15514 17587
rect 15548 17553 15554 17587
rect 15508 17515 15554 17553
rect 15508 17481 15514 17515
rect 15548 17481 15554 17515
rect 15508 17443 15554 17481
rect 15508 17409 15514 17443
rect 15548 17409 15554 17443
rect 15872 17584 15880 17601
rect 15914 17610 16980 17618
rect 15914 17602 15974 17610
rect 15914 17601 15934 17602
rect 15914 17584 15922 17601
rect 15872 17546 15922 17584
rect 15872 17512 15880 17546
rect 15914 17512 15922 17546
rect 15872 17474 15922 17512
rect 15872 17440 15880 17474
rect 15914 17440 15922 17474
rect 15872 17427 15922 17440
rect 16720 17505 16980 17610
rect 17406 17703 17456 17720
rect 17406 17669 17414 17703
rect 17448 17669 17456 17703
rect 17406 17631 17456 17669
rect 17406 17597 17414 17631
rect 17448 17597 17456 17631
rect 17406 17559 17456 17597
rect 17406 17525 17414 17559
rect 17448 17525 17456 17559
rect 17406 17512 17456 17525
rect 15508 17371 15554 17409
rect 15508 17337 15514 17371
rect 15548 17337 15554 17371
rect 15508 17299 15554 17337
rect 16720 17325 16765 17505
rect 16945 17325 16980 17505
rect 15508 17265 15514 17299
rect 15548 17265 15554 17299
rect 15508 17227 15554 17265
rect 15508 17193 15514 17227
rect 15548 17193 15554 17227
rect 15508 17155 15554 17193
rect 15508 17121 15514 17155
rect 15548 17121 15554 17155
rect 15508 17083 15554 17121
rect 15508 17049 15514 17083
rect 15548 17049 15554 17083
rect 15508 17011 15554 17049
rect 15508 16977 15514 17011
rect 15548 16977 15554 17011
rect 15872 17303 15922 17317
rect 15872 17269 15880 17303
rect 15914 17269 15922 17303
rect 15872 17231 15922 17269
rect 15872 17197 15880 17231
rect 15914 17197 15922 17231
rect 15872 17159 15922 17197
rect 15872 17125 15880 17159
rect 15914 17125 15922 17159
rect 16264 17304 16314 17318
rect 16264 17270 16272 17304
rect 16306 17270 16314 17304
rect 16720 17270 16980 17325
rect 16264 17232 16314 17270
rect 16264 17198 16272 17232
rect 16306 17198 16314 17232
rect 16264 17160 16314 17198
rect 16264 17141 16272 17160
rect 15872 17087 15922 17125
rect 15872 17053 15880 17087
rect 15914 17053 15922 17087
rect 15872 17015 15922 17053
rect 15872 16984 15880 17015
rect 15508 16934 15554 16977
rect 15816 16981 15880 16984
rect 15914 16984 15922 17015
rect 16249 17126 16272 17141
rect 16306 17141 16314 17160
rect 16306 17126 18052 17141
rect 16249 17088 18052 17126
rect 16249 17054 16272 17088
rect 16306 17054 18052 17088
rect 16249 17016 18052 17054
rect 15914 16981 15976 16984
rect 15816 16943 15976 16981
rect 14596 16401 14756 16909
rect 15816 16909 15880 16943
rect 15914 16909 15976 16943
rect 14596 16367 14623 16401
rect 14657 16367 14695 16401
rect 14729 16367 14756 16401
rect 14596 16314 14756 16367
rect 15016 16899 15126 16904
rect 15016 16896 15130 16899
rect 15016 16862 15060 16896
rect 15094 16862 15130 16896
rect 15016 16474 15130 16862
rect 15444 16896 15533 16905
rect 15444 16862 15470 16896
rect 15504 16862 15533 16896
rect 15444 16687 15533 16862
rect 15444 16635 15459 16687
rect 15511 16635 15533 16687
rect 15444 16623 15533 16635
rect 15444 16571 15459 16623
rect 15511 16571 15533 16623
rect 15444 16554 15533 16571
rect 15016 16422 15045 16474
rect 15097 16422 15130 16474
rect 15016 16410 15130 16422
rect 15016 16358 15045 16410
rect 15097 16358 15130 16410
rect 15016 16346 15130 16358
rect 13516 16279 14484 16310
rect 15016 16294 15045 16346
rect 15097 16294 15130 16346
rect 15816 16401 15976 16909
rect 16249 16982 16272 17016
rect 16306 16982 18052 17016
rect 16249 16944 18052 16982
rect 16249 16910 16272 16944
rect 16306 16910 18052 16944
rect 16249 16884 18052 16910
rect 15816 16367 15838 16401
rect 15872 16367 15910 16401
rect 15944 16367 15976 16401
rect 15816 16308 15976 16367
rect 15016 16274 15130 16294
rect 13000 16104 16242 16224
rect 13572 15536 13692 16104
rect 14742 16000 14842 16014
rect 14742 15984 14766 16000
rect 14552 15976 14766 15984
rect 14818 15984 14842 16000
rect 14818 15976 15192 15984
rect 14552 15942 14566 15976
rect 14600 15942 14758 15976
rect 14818 15948 14950 15976
rect 14792 15942 14950 15948
rect 14984 15942 15142 15976
rect 15176 15942 15192 15976
rect 14552 15934 15192 15942
rect 16122 15944 16242 16104
rect 17212 16024 17292 16044
rect 17212 15990 17236 16024
rect 17270 15990 17292 16024
rect 17212 15984 17292 15990
rect 16122 15910 16166 15944
rect 16200 15910 16242 15944
rect 13572 15502 13616 15536
rect 13650 15502 13692 15536
rect 13572 15494 13692 15502
rect 14416 15857 14462 15904
rect 14416 15823 14422 15857
rect 14456 15823 14462 15857
rect 14416 15785 14462 15823
rect 14416 15751 14422 15785
rect 14456 15751 14462 15785
rect 14493 15870 14563 15904
rect 14493 15818 14502 15870
rect 14554 15818 14563 15870
rect 14493 15785 14563 15818
rect 14493 15784 14518 15785
rect 14416 15713 14462 15751
rect 14416 15679 14422 15713
rect 14456 15679 14462 15713
rect 14416 15641 14462 15679
rect 14416 15607 14422 15641
rect 14456 15607 14462 15641
rect 14416 15569 14462 15607
rect 14416 15535 14422 15569
rect 14456 15535 14462 15569
rect 14416 15497 14462 15535
rect 13566 15452 13612 15464
rect 13507 15437 13612 15452
rect 13507 15385 13528 15437
rect 13580 15421 13612 15437
rect 13606 15387 13612 15421
rect 13580 15385 13612 15387
rect 13507 15373 13612 15385
rect 13507 15321 13528 15373
rect 13580 15349 13612 15373
rect 13507 15315 13572 15321
rect 13606 15315 13612 15349
rect 13507 15307 13612 15315
rect 13566 15277 13612 15307
rect 13566 15243 13572 15277
rect 13606 15243 13612 15277
rect 13566 15205 13612 15243
rect 13566 15171 13572 15205
rect 13606 15171 13612 15205
rect 13566 15133 13612 15171
rect 13566 15099 13572 15133
rect 13606 15099 13612 15133
rect 13566 15061 13612 15099
rect 13566 15027 13572 15061
rect 13606 15027 13612 15061
rect 13566 14989 13612 15027
rect 13566 14955 13572 14989
rect 13606 14955 13612 14989
rect 13566 14917 13612 14955
rect 13566 14883 13572 14917
rect 13606 14883 13612 14917
rect 13566 14845 13612 14883
rect 13566 14811 13572 14845
rect 13606 14811 13612 14845
rect 13566 14773 13612 14811
rect 13566 14739 13572 14773
rect 13606 14739 13612 14773
rect 13566 14701 13612 14739
rect 13566 14667 13572 14701
rect 13606 14667 13612 14701
rect 13566 14629 13612 14667
rect 13566 14595 13572 14629
rect 13606 14595 13612 14629
rect 13566 14557 13612 14595
rect 13566 14523 13572 14557
rect 13606 14523 13612 14557
rect 13566 14485 13612 14523
rect 13566 14451 13572 14485
rect 13606 14451 13612 14485
rect 13566 14413 13612 14451
rect 13566 14379 13572 14413
rect 13606 14379 13612 14413
rect 13566 14341 13612 14379
rect 13566 14307 13572 14341
rect 13606 14307 13612 14341
rect 13566 14269 13612 14307
rect 13566 14235 13572 14269
rect 13606 14235 13612 14269
rect 13566 14197 13612 14235
rect 13566 14163 13572 14197
rect 13606 14163 13612 14197
rect 13566 14125 13612 14163
rect 13566 14091 13572 14125
rect 13606 14091 13612 14125
rect 13566 14053 13612 14091
rect 13566 14020 13572 14053
rect 13480 14019 13572 14020
rect 13606 14019 13612 14053
rect 13480 13981 13612 14019
rect 13480 13947 13572 13981
rect 13606 13947 13612 13981
rect 13480 13904 13612 13947
rect 13654 15421 13700 15464
rect 13654 15387 13660 15421
rect 13694 15387 13700 15421
rect 13654 15349 13700 15387
rect 13654 15315 13660 15349
rect 13694 15315 13700 15349
rect 13654 15277 13700 15315
rect 13654 15243 13660 15277
rect 13694 15243 13700 15277
rect 13654 15205 13700 15243
rect 13654 15171 13660 15205
rect 13694 15171 13700 15205
rect 13654 15133 13700 15171
rect 13654 15099 13660 15133
rect 13694 15099 13700 15133
rect 13654 15061 13700 15099
rect 13654 15027 13660 15061
rect 13694 15027 13700 15061
rect 13654 14989 13700 15027
rect 13654 14955 13660 14989
rect 13694 14955 13700 14989
rect 13654 14917 13700 14955
rect 13654 14883 13660 14917
rect 13694 14883 13700 14917
rect 13654 14845 13700 14883
rect 13654 14811 13660 14845
rect 13694 14811 13700 14845
rect 13654 14773 13700 14811
rect 13654 14739 13660 14773
rect 13694 14739 13700 14773
rect 13654 14701 13700 14739
rect 13654 14667 13660 14701
rect 13694 14667 13700 14701
rect 13654 14629 13700 14667
rect 13654 14595 13660 14629
rect 13694 14595 13700 14629
rect 13654 14557 13700 14595
rect 13654 14523 13660 14557
rect 13694 14523 13700 14557
rect 13654 14485 13700 14523
rect 13654 14451 13660 14485
rect 13694 14451 13700 14485
rect 13654 14413 13700 14451
rect 13654 14379 13660 14413
rect 13694 14379 13700 14413
rect 13654 14341 13700 14379
rect 13654 14307 13660 14341
rect 13694 14307 13700 14341
rect 13654 14269 13700 14307
rect 13654 14235 13660 14269
rect 13694 14235 13700 14269
rect 13654 14197 13700 14235
rect 13654 14163 13660 14197
rect 13694 14163 13700 14197
rect 13654 14125 13700 14163
rect 13654 14091 13660 14125
rect 13694 14091 13700 14125
rect 13654 14053 13700 14091
rect 13654 14019 13660 14053
rect 13694 14019 13700 14053
rect 14416 15463 14422 15497
rect 14456 15463 14462 15497
rect 14416 15425 14462 15463
rect 14416 15391 14422 15425
rect 14456 15391 14462 15425
rect 14416 15353 14462 15391
rect 14416 15319 14422 15353
rect 14456 15319 14462 15353
rect 14416 15281 14462 15319
rect 14416 15247 14422 15281
rect 14456 15247 14462 15281
rect 14416 15209 14462 15247
rect 14416 15175 14422 15209
rect 14456 15175 14462 15209
rect 14416 15137 14462 15175
rect 14416 15103 14422 15137
rect 14456 15103 14462 15137
rect 14416 15065 14462 15103
rect 14416 15031 14422 15065
rect 14456 15031 14462 15065
rect 14416 14993 14462 15031
rect 14416 14959 14422 14993
rect 14456 14959 14462 14993
rect 14416 14921 14462 14959
rect 14416 14887 14422 14921
rect 14456 14887 14462 14921
rect 14416 14849 14462 14887
rect 14416 14815 14422 14849
rect 14456 14815 14462 14849
rect 14416 14777 14462 14815
rect 14416 14743 14422 14777
rect 14456 14743 14462 14777
rect 14416 14705 14462 14743
rect 14416 14671 14422 14705
rect 14456 14671 14462 14705
rect 14416 14633 14462 14671
rect 14416 14599 14422 14633
rect 14456 14599 14462 14633
rect 14416 14561 14462 14599
rect 14416 14527 14422 14561
rect 14456 14527 14462 14561
rect 14416 14489 14462 14527
rect 14416 14455 14422 14489
rect 14456 14455 14462 14489
rect 14416 14417 14462 14455
rect 14416 14383 14422 14417
rect 14456 14383 14462 14417
rect 14416 14345 14462 14383
rect 14416 14311 14422 14345
rect 14456 14311 14462 14345
rect 14416 14273 14462 14311
rect 14416 14239 14422 14273
rect 14456 14239 14462 14273
rect 14416 14201 14462 14239
rect 14416 14167 14422 14201
rect 14456 14167 14462 14201
rect 14416 14129 14462 14167
rect 14416 14095 14422 14129
rect 14456 14095 14462 14129
rect 14416 14057 14462 14095
rect 14416 14034 14422 14057
rect 13654 13981 13700 14019
rect 13654 13947 13660 13981
rect 13694 13947 13700 13981
rect 13654 13904 13700 13947
rect 14413 14023 14422 14034
rect 14456 14034 14462 14057
rect 14512 15751 14518 15784
rect 14552 15784 14563 15785
rect 14608 15857 14654 15904
rect 14608 15823 14614 15857
rect 14648 15823 14654 15857
rect 14608 15785 14654 15823
rect 14552 15751 14558 15784
rect 14512 15713 14558 15751
rect 14512 15679 14518 15713
rect 14552 15679 14558 15713
rect 14512 15641 14558 15679
rect 14512 15607 14518 15641
rect 14552 15607 14558 15641
rect 14512 15569 14558 15607
rect 14512 15535 14518 15569
rect 14552 15535 14558 15569
rect 14512 15497 14558 15535
rect 14512 15463 14518 15497
rect 14552 15463 14558 15497
rect 14512 15425 14558 15463
rect 14512 15391 14518 15425
rect 14552 15391 14558 15425
rect 14512 15353 14558 15391
rect 14512 15319 14518 15353
rect 14552 15319 14558 15353
rect 14512 15281 14558 15319
rect 14512 15247 14518 15281
rect 14552 15247 14558 15281
rect 14512 15209 14558 15247
rect 14512 15175 14518 15209
rect 14552 15175 14558 15209
rect 14512 15137 14558 15175
rect 14512 15103 14518 15137
rect 14552 15103 14558 15137
rect 14512 15065 14558 15103
rect 14512 15031 14518 15065
rect 14552 15031 14558 15065
rect 14512 14993 14558 15031
rect 14512 14959 14518 14993
rect 14552 14959 14558 14993
rect 14512 14921 14558 14959
rect 14512 14887 14518 14921
rect 14552 14887 14558 14921
rect 14512 14849 14558 14887
rect 14512 14815 14518 14849
rect 14552 14815 14558 14849
rect 14512 14777 14558 14815
rect 14512 14743 14518 14777
rect 14552 14743 14558 14777
rect 14512 14705 14558 14743
rect 14512 14671 14518 14705
rect 14552 14671 14558 14705
rect 14512 14633 14558 14671
rect 14512 14599 14518 14633
rect 14552 14599 14558 14633
rect 14512 14561 14558 14599
rect 14512 14527 14518 14561
rect 14552 14527 14558 14561
rect 14512 14489 14558 14527
rect 14512 14455 14518 14489
rect 14552 14455 14558 14489
rect 14512 14417 14558 14455
rect 14512 14383 14518 14417
rect 14552 14383 14558 14417
rect 14512 14345 14558 14383
rect 14512 14311 14518 14345
rect 14552 14311 14558 14345
rect 14512 14273 14558 14311
rect 14512 14239 14518 14273
rect 14552 14239 14558 14273
rect 14512 14201 14558 14239
rect 14512 14167 14518 14201
rect 14552 14167 14558 14201
rect 14512 14129 14558 14167
rect 14512 14095 14518 14129
rect 14552 14095 14558 14129
rect 14512 14057 14558 14095
rect 14456 14023 14483 14034
rect 14413 14000 14483 14023
rect 14413 13948 14422 14000
rect 14474 13948 14483 14000
rect 14413 13914 14483 13948
rect 14512 14023 14518 14057
rect 14552 14023 14558 14057
rect 14608 15751 14614 15785
rect 14648 15751 14654 15785
rect 14693 15870 14763 15904
rect 14693 15818 14702 15870
rect 14754 15818 14763 15870
rect 14693 15785 14763 15818
rect 14693 15784 14710 15785
rect 14608 15713 14654 15751
rect 14608 15679 14614 15713
rect 14648 15679 14654 15713
rect 14608 15641 14654 15679
rect 14608 15607 14614 15641
rect 14648 15607 14654 15641
rect 14608 15569 14654 15607
rect 14608 15535 14614 15569
rect 14648 15535 14654 15569
rect 14608 15497 14654 15535
rect 14608 15463 14614 15497
rect 14648 15463 14654 15497
rect 14608 15425 14654 15463
rect 14608 15391 14614 15425
rect 14648 15391 14654 15425
rect 14608 15353 14654 15391
rect 14608 15319 14614 15353
rect 14648 15319 14654 15353
rect 14608 15281 14654 15319
rect 14608 15247 14614 15281
rect 14648 15247 14654 15281
rect 14608 15209 14654 15247
rect 14608 15175 14614 15209
rect 14648 15175 14654 15209
rect 14608 15137 14654 15175
rect 14608 15103 14614 15137
rect 14648 15103 14654 15137
rect 14608 15065 14654 15103
rect 14608 15031 14614 15065
rect 14648 15031 14654 15065
rect 14608 14993 14654 15031
rect 14608 14959 14614 14993
rect 14648 14959 14654 14993
rect 14608 14921 14654 14959
rect 14608 14887 14614 14921
rect 14648 14887 14654 14921
rect 14608 14849 14654 14887
rect 14608 14815 14614 14849
rect 14648 14815 14654 14849
rect 14608 14777 14654 14815
rect 14608 14743 14614 14777
rect 14648 14743 14654 14777
rect 14608 14705 14654 14743
rect 14608 14671 14614 14705
rect 14648 14671 14654 14705
rect 14608 14633 14654 14671
rect 14608 14599 14614 14633
rect 14648 14599 14654 14633
rect 14608 14561 14654 14599
rect 14608 14527 14614 14561
rect 14648 14527 14654 14561
rect 14608 14489 14654 14527
rect 14608 14455 14614 14489
rect 14648 14455 14654 14489
rect 14608 14417 14654 14455
rect 14608 14383 14614 14417
rect 14648 14383 14654 14417
rect 14608 14345 14654 14383
rect 14608 14311 14614 14345
rect 14648 14311 14654 14345
rect 14608 14273 14654 14311
rect 14608 14239 14614 14273
rect 14648 14239 14654 14273
rect 14608 14201 14654 14239
rect 14608 14167 14614 14201
rect 14648 14167 14654 14201
rect 14608 14129 14654 14167
rect 14608 14095 14614 14129
rect 14648 14095 14654 14129
rect 14608 14057 14654 14095
rect 14608 14034 14614 14057
rect 14512 13985 14558 14023
rect 14512 13951 14518 13985
rect 14552 13951 14558 13985
rect 14416 13904 14462 13914
rect 14512 13904 14558 13951
rect 14593 14023 14614 14034
rect 14648 14034 14654 14057
rect 14704 15751 14710 15784
rect 14744 15784 14763 15785
rect 14800 15857 14846 15904
rect 14800 15823 14806 15857
rect 14840 15823 14846 15857
rect 14800 15785 14846 15823
rect 14744 15751 14750 15784
rect 14704 15713 14750 15751
rect 14704 15679 14710 15713
rect 14744 15679 14750 15713
rect 14704 15641 14750 15679
rect 14704 15607 14710 15641
rect 14744 15607 14750 15641
rect 14704 15569 14750 15607
rect 14704 15535 14710 15569
rect 14744 15535 14750 15569
rect 14704 15497 14750 15535
rect 14704 15463 14710 15497
rect 14744 15463 14750 15497
rect 14704 15425 14750 15463
rect 14704 15391 14710 15425
rect 14744 15391 14750 15425
rect 14704 15353 14750 15391
rect 14704 15319 14710 15353
rect 14744 15319 14750 15353
rect 14704 15281 14750 15319
rect 14704 15247 14710 15281
rect 14744 15247 14750 15281
rect 14704 15209 14750 15247
rect 14704 15175 14710 15209
rect 14744 15175 14750 15209
rect 14704 15137 14750 15175
rect 14704 15103 14710 15137
rect 14744 15103 14750 15137
rect 14704 15065 14750 15103
rect 14704 15031 14710 15065
rect 14744 15031 14750 15065
rect 14704 14993 14750 15031
rect 14704 14959 14710 14993
rect 14744 14959 14750 14993
rect 14704 14921 14750 14959
rect 14704 14887 14710 14921
rect 14744 14887 14750 14921
rect 14704 14849 14750 14887
rect 14704 14815 14710 14849
rect 14744 14815 14750 14849
rect 14704 14777 14750 14815
rect 14704 14743 14710 14777
rect 14744 14743 14750 14777
rect 14704 14705 14750 14743
rect 14704 14671 14710 14705
rect 14744 14671 14750 14705
rect 14704 14633 14750 14671
rect 14704 14599 14710 14633
rect 14744 14599 14750 14633
rect 14704 14561 14750 14599
rect 14704 14527 14710 14561
rect 14744 14527 14750 14561
rect 14704 14489 14750 14527
rect 14704 14455 14710 14489
rect 14744 14455 14750 14489
rect 14704 14417 14750 14455
rect 14704 14383 14710 14417
rect 14744 14383 14750 14417
rect 14704 14345 14750 14383
rect 14704 14311 14710 14345
rect 14744 14311 14750 14345
rect 14704 14273 14750 14311
rect 14704 14239 14710 14273
rect 14744 14239 14750 14273
rect 14704 14201 14750 14239
rect 14704 14167 14710 14201
rect 14744 14167 14750 14201
rect 14704 14129 14750 14167
rect 14704 14095 14710 14129
rect 14744 14095 14750 14129
rect 14704 14057 14750 14095
rect 14648 14023 14663 14034
rect 14593 14000 14663 14023
rect 14593 13948 14602 14000
rect 14654 13948 14663 14000
rect 14593 13914 14663 13948
rect 14704 14023 14710 14057
rect 14744 14023 14750 14057
rect 14800 15751 14806 15785
rect 14840 15751 14846 15785
rect 14883 15870 14953 15904
rect 14883 15818 14892 15870
rect 14944 15818 14953 15870
rect 14883 15785 14953 15818
rect 14883 15784 14902 15785
rect 14800 15713 14846 15751
rect 14800 15679 14806 15713
rect 14840 15679 14846 15713
rect 14800 15641 14846 15679
rect 14800 15607 14806 15641
rect 14840 15607 14846 15641
rect 14800 15569 14846 15607
rect 14800 15535 14806 15569
rect 14840 15535 14846 15569
rect 14800 15497 14846 15535
rect 14800 15463 14806 15497
rect 14840 15463 14846 15497
rect 14800 15425 14846 15463
rect 14800 15391 14806 15425
rect 14840 15391 14846 15425
rect 14800 15353 14846 15391
rect 14800 15319 14806 15353
rect 14840 15319 14846 15353
rect 14800 15281 14846 15319
rect 14800 15247 14806 15281
rect 14840 15247 14846 15281
rect 14800 15209 14846 15247
rect 14800 15175 14806 15209
rect 14840 15175 14846 15209
rect 14800 15137 14846 15175
rect 14800 15103 14806 15137
rect 14840 15103 14846 15137
rect 14800 15065 14846 15103
rect 14800 15031 14806 15065
rect 14840 15031 14846 15065
rect 14800 14993 14846 15031
rect 14800 14959 14806 14993
rect 14840 14959 14846 14993
rect 14800 14921 14846 14959
rect 14800 14887 14806 14921
rect 14840 14887 14846 14921
rect 14800 14849 14846 14887
rect 14800 14815 14806 14849
rect 14840 14815 14846 14849
rect 14800 14777 14846 14815
rect 14800 14743 14806 14777
rect 14840 14743 14846 14777
rect 14800 14705 14846 14743
rect 14800 14671 14806 14705
rect 14840 14671 14846 14705
rect 14800 14633 14846 14671
rect 14800 14599 14806 14633
rect 14840 14599 14846 14633
rect 14800 14561 14846 14599
rect 14800 14527 14806 14561
rect 14840 14527 14846 14561
rect 14800 14489 14846 14527
rect 14800 14455 14806 14489
rect 14840 14455 14846 14489
rect 14800 14417 14846 14455
rect 14800 14383 14806 14417
rect 14840 14383 14846 14417
rect 14800 14345 14846 14383
rect 14800 14311 14806 14345
rect 14840 14311 14846 14345
rect 14800 14273 14846 14311
rect 14800 14239 14806 14273
rect 14840 14239 14846 14273
rect 14800 14201 14846 14239
rect 14800 14167 14806 14201
rect 14840 14167 14846 14201
rect 14800 14129 14846 14167
rect 14800 14095 14806 14129
rect 14840 14095 14846 14129
rect 14800 14057 14846 14095
rect 14800 14034 14806 14057
rect 14704 13985 14750 14023
rect 14704 13951 14710 13985
rect 14744 13951 14750 13985
rect 14608 13904 14654 13914
rect 14704 13904 14750 13951
rect 14783 14023 14806 14034
rect 14840 14034 14846 14057
rect 14896 15751 14902 15784
rect 14936 15784 14953 15785
rect 14992 15857 15038 15904
rect 14992 15823 14998 15857
rect 15032 15823 15038 15857
rect 14992 15785 15038 15823
rect 14936 15751 14942 15784
rect 14896 15713 14942 15751
rect 14896 15679 14902 15713
rect 14936 15679 14942 15713
rect 14896 15641 14942 15679
rect 14896 15607 14902 15641
rect 14936 15607 14942 15641
rect 14896 15569 14942 15607
rect 14896 15535 14902 15569
rect 14936 15535 14942 15569
rect 14896 15497 14942 15535
rect 14896 15463 14902 15497
rect 14936 15463 14942 15497
rect 14896 15425 14942 15463
rect 14896 15391 14902 15425
rect 14936 15391 14942 15425
rect 14896 15353 14942 15391
rect 14896 15319 14902 15353
rect 14936 15319 14942 15353
rect 14896 15281 14942 15319
rect 14896 15247 14902 15281
rect 14936 15247 14942 15281
rect 14896 15209 14942 15247
rect 14896 15175 14902 15209
rect 14936 15175 14942 15209
rect 14896 15137 14942 15175
rect 14896 15103 14902 15137
rect 14936 15103 14942 15137
rect 14896 15065 14942 15103
rect 14896 15031 14902 15065
rect 14936 15031 14942 15065
rect 14896 14993 14942 15031
rect 14896 14959 14902 14993
rect 14936 14959 14942 14993
rect 14896 14921 14942 14959
rect 14896 14887 14902 14921
rect 14936 14887 14942 14921
rect 14896 14849 14942 14887
rect 14896 14815 14902 14849
rect 14936 14815 14942 14849
rect 14896 14777 14942 14815
rect 14896 14743 14902 14777
rect 14936 14743 14942 14777
rect 14896 14705 14942 14743
rect 14896 14671 14902 14705
rect 14936 14671 14942 14705
rect 14896 14633 14942 14671
rect 14896 14599 14902 14633
rect 14936 14599 14942 14633
rect 14896 14561 14942 14599
rect 14896 14527 14902 14561
rect 14936 14527 14942 14561
rect 14896 14489 14942 14527
rect 14896 14455 14902 14489
rect 14936 14455 14942 14489
rect 14896 14417 14942 14455
rect 14896 14383 14902 14417
rect 14936 14383 14942 14417
rect 14896 14345 14942 14383
rect 14896 14311 14902 14345
rect 14936 14311 14942 14345
rect 14896 14273 14942 14311
rect 14896 14239 14902 14273
rect 14936 14239 14942 14273
rect 14896 14201 14942 14239
rect 14896 14167 14902 14201
rect 14936 14167 14942 14201
rect 14896 14129 14942 14167
rect 14896 14095 14902 14129
rect 14936 14095 14942 14129
rect 14896 14057 14942 14095
rect 14840 14023 14853 14034
rect 14783 14000 14853 14023
rect 14783 13948 14792 14000
rect 14844 13948 14853 14000
rect 14783 13914 14853 13948
rect 14896 14023 14902 14057
rect 14936 14023 14942 14057
rect 14992 15751 14998 15785
rect 15032 15751 15038 15785
rect 15073 15870 15143 15904
rect 15073 15818 15082 15870
rect 15134 15818 15143 15870
rect 15073 15785 15143 15818
rect 15073 15784 15094 15785
rect 14992 15713 15038 15751
rect 14992 15679 14998 15713
rect 15032 15679 15038 15713
rect 14992 15641 15038 15679
rect 14992 15607 14998 15641
rect 15032 15607 15038 15641
rect 14992 15569 15038 15607
rect 14992 15535 14998 15569
rect 15032 15535 15038 15569
rect 14992 15497 15038 15535
rect 14992 15463 14998 15497
rect 15032 15463 15038 15497
rect 14992 15425 15038 15463
rect 14992 15391 14998 15425
rect 15032 15391 15038 15425
rect 14992 15353 15038 15391
rect 14992 15319 14998 15353
rect 15032 15319 15038 15353
rect 14992 15281 15038 15319
rect 14992 15247 14998 15281
rect 15032 15247 15038 15281
rect 14992 15209 15038 15247
rect 14992 15175 14998 15209
rect 15032 15175 15038 15209
rect 14992 15137 15038 15175
rect 14992 15103 14998 15137
rect 15032 15103 15038 15137
rect 14992 15065 15038 15103
rect 14992 15031 14998 15065
rect 15032 15031 15038 15065
rect 14992 14993 15038 15031
rect 14992 14959 14998 14993
rect 15032 14959 15038 14993
rect 14992 14921 15038 14959
rect 14992 14887 14998 14921
rect 15032 14887 15038 14921
rect 14992 14849 15038 14887
rect 14992 14815 14998 14849
rect 15032 14815 15038 14849
rect 14992 14777 15038 14815
rect 14992 14743 14998 14777
rect 15032 14743 15038 14777
rect 14992 14705 15038 14743
rect 14992 14671 14998 14705
rect 15032 14671 15038 14705
rect 14992 14633 15038 14671
rect 14992 14599 14998 14633
rect 15032 14599 15038 14633
rect 14992 14561 15038 14599
rect 14992 14527 14998 14561
rect 15032 14527 15038 14561
rect 14992 14489 15038 14527
rect 14992 14455 14998 14489
rect 15032 14455 15038 14489
rect 14992 14417 15038 14455
rect 14992 14383 14998 14417
rect 15032 14383 15038 14417
rect 14992 14345 15038 14383
rect 14992 14311 14998 14345
rect 15032 14311 15038 14345
rect 14992 14273 15038 14311
rect 14992 14239 14998 14273
rect 15032 14239 15038 14273
rect 14992 14201 15038 14239
rect 14992 14167 14998 14201
rect 15032 14167 15038 14201
rect 14992 14129 15038 14167
rect 14992 14095 14998 14129
rect 15032 14095 15038 14129
rect 14992 14057 15038 14095
rect 14992 14034 14998 14057
rect 14896 13985 14942 14023
rect 14896 13951 14902 13985
rect 14936 13951 14942 13985
rect 14800 13904 14846 13914
rect 14896 13904 14942 13951
rect 14973 14023 14998 14034
rect 15032 14034 15038 14057
rect 15088 15751 15094 15784
rect 15128 15784 15143 15785
rect 15184 15857 15230 15904
rect 15184 15823 15190 15857
rect 15224 15823 15230 15857
rect 15184 15785 15230 15823
rect 15128 15751 15134 15784
rect 15088 15713 15134 15751
rect 15088 15679 15094 15713
rect 15128 15679 15134 15713
rect 15088 15641 15134 15679
rect 15088 15607 15094 15641
rect 15128 15607 15134 15641
rect 15088 15569 15134 15607
rect 15088 15535 15094 15569
rect 15128 15535 15134 15569
rect 15088 15497 15134 15535
rect 15088 15463 15094 15497
rect 15128 15463 15134 15497
rect 15088 15425 15134 15463
rect 15088 15391 15094 15425
rect 15128 15391 15134 15425
rect 15088 15353 15134 15391
rect 15088 15319 15094 15353
rect 15128 15319 15134 15353
rect 15088 15281 15134 15319
rect 15088 15247 15094 15281
rect 15128 15247 15134 15281
rect 15088 15209 15134 15247
rect 15088 15175 15094 15209
rect 15128 15175 15134 15209
rect 15088 15137 15134 15175
rect 15088 15103 15094 15137
rect 15128 15103 15134 15137
rect 15088 15065 15134 15103
rect 15088 15031 15094 15065
rect 15128 15031 15134 15065
rect 15088 14993 15134 15031
rect 15088 14959 15094 14993
rect 15128 14959 15134 14993
rect 15088 14921 15134 14959
rect 15088 14887 15094 14921
rect 15128 14887 15134 14921
rect 15088 14849 15134 14887
rect 15088 14815 15094 14849
rect 15128 14815 15134 14849
rect 15088 14777 15134 14815
rect 15088 14743 15094 14777
rect 15128 14743 15134 14777
rect 15088 14705 15134 14743
rect 15088 14671 15094 14705
rect 15128 14671 15134 14705
rect 15088 14633 15134 14671
rect 15088 14599 15094 14633
rect 15128 14599 15134 14633
rect 15088 14561 15134 14599
rect 15088 14527 15094 14561
rect 15128 14527 15134 14561
rect 15088 14489 15134 14527
rect 15088 14455 15094 14489
rect 15128 14455 15134 14489
rect 15088 14417 15134 14455
rect 15088 14383 15094 14417
rect 15128 14383 15134 14417
rect 15088 14345 15134 14383
rect 15088 14311 15094 14345
rect 15128 14311 15134 14345
rect 15088 14273 15134 14311
rect 15088 14239 15094 14273
rect 15128 14239 15134 14273
rect 15088 14201 15134 14239
rect 15088 14167 15094 14201
rect 15128 14167 15134 14201
rect 15088 14129 15134 14167
rect 15088 14095 15094 14129
rect 15128 14095 15134 14129
rect 15088 14057 15134 14095
rect 15032 14023 15043 14034
rect 14973 14000 15043 14023
rect 14973 13948 14982 14000
rect 15034 13948 15043 14000
rect 14973 13914 15043 13948
rect 15088 14023 15094 14057
rect 15128 14023 15134 14057
rect 15184 15751 15190 15785
rect 15224 15751 15230 15785
rect 15184 15713 15230 15751
rect 15184 15679 15190 15713
rect 15224 15679 15230 15713
rect 15184 15641 15230 15679
rect 15184 15607 15190 15641
rect 15224 15607 15230 15641
rect 15184 15569 15230 15607
rect 15184 15535 15190 15569
rect 15224 15535 15230 15569
rect 15184 15497 15230 15535
rect 16122 15872 16242 15910
rect 16122 15838 16166 15872
rect 16200 15838 16242 15872
rect 16122 15800 16242 15838
rect 16122 15766 16166 15800
rect 16200 15766 16242 15800
rect 16122 15728 16242 15766
rect 16122 15694 16166 15728
rect 16200 15694 16242 15728
rect 16122 15656 16242 15694
rect 16122 15622 16166 15656
rect 16200 15622 16242 15656
rect 16122 15584 16242 15622
rect 16122 15550 16166 15584
rect 16200 15550 16242 15584
rect 16122 15524 16242 15550
rect 17086 15896 17132 15943
rect 17086 15862 17092 15896
rect 17126 15862 17132 15896
rect 17086 15824 17132 15862
rect 17173 15910 17243 15944
rect 17173 15858 17182 15910
rect 17234 15858 17243 15910
rect 17173 15824 17243 15858
rect 17278 15896 17324 15943
rect 17278 15862 17284 15896
rect 17318 15862 17324 15896
rect 17278 15824 17324 15862
rect 17363 15910 17433 15944
rect 17363 15858 17372 15910
rect 17424 15858 17433 15910
rect 17363 15824 17433 15858
rect 17086 15790 17092 15824
rect 17126 15790 17132 15824
rect 17086 15752 17132 15790
rect 17086 15718 17092 15752
rect 17126 15718 17132 15752
rect 17086 15680 17132 15718
rect 17086 15646 17092 15680
rect 17126 15646 17132 15680
rect 17086 15608 17132 15646
rect 17086 15574 17092 15608
rect 17126 15574 17132 15608
rect 17086 15536 17132 15574
rect 15184 15463 15190 15497
rect 15224 15463 15230 15497
rect 15184 15425 15230 15463
rect 15184 15391 15190 15425
rect 15224 15391 15230 15425
rect 15184 15353 15230 15391
rect 15184 15319 15190 15353
rect 15224 15319 15230 15353
rect 15184 15281 15230 15319
rect 15184 15247 15190 15281
rect 15224 15247 15230 15281
rect 15184 15209 15230 15247
rect 15184 15175 15190 15209
rect 15224 15175 15230 15209
rect 15184 15137 15230 15175
rect 15184 15103 15190 15137
rect 15224 15103 15230 15137
rect 15184 15065 15230 15103
rect 15184 15031 15190 15065
rect 15224 15031 15230 15065
rect 15184 14993 15230 15031
rect 15184 14959 15190 14993
rect 15224 14959 15230 14993
rect 15184 14921 15230 14959
rect 15184 14887 15190 14921
rect 15224 14887 15230 14921
rect 15184 14849 15230 14887
rect 15184 14815 15190 14849
rect 15224 14815 15230 14849
rect 15184 14777 15230 14815
rect 15184 14743 15190 14777
rect 15224 14743 15230 14777
rect 15184 14705 15230 14743
rect 15184 14671 15190 14705
rect 15224 14671 15230 14705
rect 15184 14633 15230 14671
rect 15184 14599 15190 14633
rect 15224 14599 15230 14633
rect 15184 14561 15230 14599
rect 15184 14527 15190 14561
rect 15224 14527 15230 14561
rect 15184 14489 15230 14527
rect 15184 14455 15190 14489
rect 15224 14455 15230 14489
rect 15184 14417 15230 14455
rect 15184 14383 15190 14417
rect 15224 14383 15230 14417
rect 15184 14345 15230 14383
rect 15184 14311 15190 14345
rect 15224 14311 15230 14345
rect 17086 15502 17092 15536
rect 17126 15502 17132 15536
rect 17086 15464 17132 15502
rect 17086 15430 17092 15464
rect 17126 15430 17132 15464
rect 17086 15392 17132 15430
rect 17086 15358 17092 15392
rect 17126 15358 17132 15392
rect 17086 15320 17132 15358
rect 17086 15286 17092 15320
rect 17126 15286 17132 15320
rect 17086 15248 17132 15286
rect 17086 15214 17092 15248
rect 17126 15214 17132 15248
rect 17086 15176 17132 15214
rect 17086 15142 17092 15176
rect 17126 15142 17132 15176
rect 17086 15104 17132 15142
rect 17086 15070 17092 15104
rect 17126 15070 17132 15104
rect 17086 15032 17132 15070
rect 17086 14998 17092 15032
rect 17126 14998 17132 15032
rect 17086 14960 17132 14998
rect 17086 14926 17092 14960
rect 17126 14926 17132 14960
rect 17086 14888 17132 14926
rect 17086 14854 17092 14888
rect 17126 14854 17132 14888
rect 17086 14816 17132 14854
rect 17086 14782 17092 14816
rect 17126 14782 17132 14816
rect 17086 14744 17132 14782
rect 17086 14710 17092 14744
rect 17126 14710 17132 14744
rect 17086 14672 17132 14710
rect 17086 14638 17092 14672
rect 17126 14638 17132 14672
rect 17086 14600 17132 14638
rect 17086 14566 17092 14600
rect 17126 14566 17132 14600
rect 17086 14528 17132 14566
rect 17086 14494 17092 14528
rect 17126 14494 17132 14528
rect 17086 14456 17132 14494
rect 17086 14422 17092 14456
rect 17126 14422 17132 14456
rect 17086 14384 17132 14422
rect 17086 14350 17092 14384
rect 17126 14350 17132 14384
rect 15184 14273 15230 14311
rect 15184 14239 15190 14273
rect 15224 14239 15230 14273
rect 15184 14201 15230 14239
rect 15184 14167 15190 14201
rect 15224 14167 15230 14201
rect 15184 14129 15230 14167
rect 15184 14095 15190 14129
rect 15224 14095 15230 14129
rect 15184 14057 15230 14095
rect 15184 14034 15190 14057
rect 15088 13985 15134 14023
rect 15088 13951 15094 13985
rect 15128 13951 15134 13985
rect 14992 13904 15038 13914
rect 15088 13904 15134 13951
rect 15163 14023 15190 14034
rect 15224 14034 15230 14057
rect 16122 14273 16242 14314
rect 16122 14239 16166 14273
rect 16200 14239 16242 14273
rect 16122 14201 16242 14239
rect 16122 14167 16166 14201
rect 16200 14167 16242 14201
rect 16122 14129 16242 14167
rect 16122 14095 16166 14129
rect 16200 14095 16242 14129
rect 16122 14057 16242 14095
rect 17086 14312 17132 14350
rect 17086 14278 17092 14312
rect 17126 14278 17132 14312
rect 17086 14240 17132 14278
rect 17086 14206 17092 14240
rect 17126 14206 17132 14240
rect 17086 14168 17132 14206
rect 17086 14134 17092 14168
rect 17126 14134 17132 14168
rect 17086 14096 17132 14134
rect 17086 14064 17092 14096
rect 15224 14023 15233 14034
rect 15163 14000 15233 14023
rect 15163 13948 15172 14000
rect 15224 13948 15233 14000
rect 15163 13914 15233 13948
rect 16122 14023 16166 14057
rect 16200 14023 16242 14057
rect 16122 13985 16242 14023
rect 16122 13951 16166 13985
rect 16200 13951 16242 13985
rect 15184 13904 15230 13914
rect 16122 13913 16242 13951
rect 17073 14062 17092 14064
rect 17126 14064 17132 14096
rect 17182 15790 17188 15824
rect 17222 15790 17228 15824
rect 17182 15752 17228 15790
rect 17182 15718 17188 15752
rect 17222 15718 17228 15752
rect 17182 15680 17228 15718
rect 17182 15646 17188 15680
rect 17222 15646 17228 15680
rect 17182 15608 17228 15646
rect 17182 15574 17188 15608
rect 17222 15574 17228 15608
rect 17182 15536 17228 15574
rect 17182 15502 17188 15536
rect 17222 15502 17228 15536
rect 17182 15464 17228 15502
rect 17182 15430 17188 15464
rect 17222 15430 17228 15464
rect 17182 15392 17228 15430
rect 17182 15358 17188 15392
rect 17222 15358 17228 15392
rect 17182 15320 17228 15358
rect 17182 15286 17188 15320
rect 17222 15286 17228 15320
rect 17182 15248 17228 15286
rect 17182 15214 17188 15248
rect 17222 15214 17228 15248
rect 17182 15176 17228 15214
rect 17182 15142 17188 15176
rect 17222 15142 17228 15176
rect 17182 15104 17228 15142
rect 17182 15070 17188 15104
rect 17222 15070 17228 15104
rect 17182 15032 17228 15070
rect 17182 14998 17188 15032
rect 17222 14998 17228 15032
rect 17182 14960 17228 14998
rect 17182 14926 17188 14960
rect 17222 14926 17228 14960
rect 17182 14888 17228 14926
rect 17182 14854 17188 14888
rect 17222 14854 17228 14888
rect 17182 14816 17228 14854
rect 17182 14782 17188 14816
rect 17222 14782 17228 14816
rect 17182 14744 17228 14782
rect 17182 14710 17188 14744
rect 17222 14710 17228 14744
rect 17182 14672 17228 14710
rect 17182 14638 17188 14672
rect 17222 14638 17228 14672
rect 17182 14600 17228 14638
rect 17182 14566 17188 14600
rect 17222 14566 17228 14600
rect 17182 14528 17228 14566
rect 17182 14494 17188 14528
rect 17222 14494 17228 14528
rect 17182 14456 17228 14494
rect 17182 14422 17188 14456
rect 17222 14422 17228 14456
rect 17182 14384 17228 14422
rect 17182 14350 17188 14384
rect 17222 14350 17228 14384
rect 17182 14312 17228 14350
rect 17182 14278 17188 14312
rect 17222 14278 17228 14312
rect 17182 14240 17228 14278
rect 17182 14206 17188 14240
rect 17222 14206 17228 14240
rect 17182 14168 17228 14206
rect 17182 14134 17188 14168
rect 17222 14134 17228 14168
rect 17182 14096 17228 14134
rect 17126 14062 17143 14064
rect 17073 14030 17143 14062
rect 17073 13978 17082 14030
rect 17134 13978 17143 14030
rect 17073 13944 17143 13978
rect 17182 14062 17188 14096
rect 17222 14062 17228 14096
rect 17278 15790 17284 15824
rect 17318 15790 17324 15824
rect 17278 15752 17324 15790
rect 17278 15718 17284 15752
rect 17318 15718 17324 15752
rect 17278 15680 17324 15718
rect 17278 15646 17284 15680
rect 17318 15646 17324 15680
rect 17278 15608 17324 15646
rect 17278 15574 17284 15608
rect 17318 15574 17324 15608
rect 17278 15536 17324 15574
rect 17278 15502 17284 15536
rect 17318 15502 17324 15536
rect 17278 15464 17324 15502
rect 17278 15430 17284 15464
rect 17318 15430 17324 15464
rect 17278 15392 17324 15430
rect 17278 15358 17284 15392
rect 17318 15358 17324 15392
rect 17278 15320 17324 15358
rect 17278 15286 17284 15320
rect 17318 15286 17324 15320
rect 17278 15248 17324 15286
rect 17278 15214 17284 15248
rect 17318 15214 17324 15248
rect 17278 15176 17324 15214
rect 17278 15142 17284 15176
rect 17318 15142 17324 15176
rect 17278 15104 17324 15142
rect 17278 15070 17284 15104
rect 17318 15070 17324 15104
rect 17278 15032 17324 15070
rect 17278 14998 17284 15032
rect 17318 14998 17324 15032
rect 17278 14960 17324 14998
rect 17278 14926 17284 14960
rect 17318 14926 17324 14960
rect 17278 14888 17324 14926
rect 17278 14854 17284 14888
rect 17318 14854 17324 14888
rect 17278 14816 17324 14854
rect 17278 14782 17284 14816
rect 17318 14782 17324 14816
rect 17278 14744 17324 14782
rect 17278 14710 17284 14744
rect 17318 14710 17324 14744
rect 17278 14672 17324 14710
rect 17278 14638 17284 14672
rect 17318 14638 17324 14672
rect 17278 14600 17324 14638
rect 17278 14566 17284 14600
rect 17318 14566 17324 14600
rect 17278 14528 17324 14566
rect 17278 14494 17284 14528
rect 17318 14494 17324 14528
rect 17278 14456 17324 14494
rect 17278 14422 17284 14456
rect 17318 14422 17324 14456
rect 17278 14384 17324 14422
rect 17278 14350 17284 14384
rect 17318 14350 17324 14384
rect 17278 14312 17324 14350
rect 17278 14278 17284 14312
rect 17318 14278 17324 14312
rect 17278 14240 17324 14278
rect 17278 14206 17284 14240
rect 17318 14206 17324 14240
rect 17278 14168 17324 14206
rect 17278 14134 17284 14168
rect 17318 14134 17324 14168
rect 17278 14096 17324 14134
rect 17278 14064 17284 14096
rect 17182 14024 17228 14062
rect 17182 13990 17188 14024
rect 17222 13990 17228 14024
rect 17086 13943 17132 13944
rect 17182 13943 17228 13990
rect 17273 14062 17284 14064
rect 17318 14064 17324 14096
rect 17374 15790 17380 15824
rect 17414 15790 17420 15824
rect 17374 15752 17420 15790
rect 17374 15718 17380 15752
rect 17414 15718 17420 15752
rect 17374 15680 17420 15718
rect 17374 15646 17380 15680
rect 17414 15646 17420 15680
rect 17374 15608 17420 15646
rect 17374 15574 17380 15608
rect 17414 15574 17420 15608
rect 17374 15536 17420 15574
rect 17374 15502 17380 15536
rect 17414 15502 17420 15536
rect 17374 15464 17420 15502
rect 17374 15430 17380 15464
rect 17414 15430 17420 15464
rect 17374 15392 17420 15430
rect 17374 15358 17380 15392
rect 17414 15358 17420 15392
rect 17374 15320 17420 15358
rect 17374 15286 17380 15320
rect 17414 15286 17420 15320
rect 17374 15248 17420 15286
rect 17374 15214 17380 15248
rect 17414 15214 17420 15248
rect 17374 15176 17420 15214
rect 17374 15142 17380 15176
rect 17414 15142 17420 15176
rect 17374 15104 17420 15142
rect 17374 15070 17380 15104
rect 17414 15070 17420 15104
rect 17374 15032 17420 15070
rect 17374 14998 17380 15032
rect 17414 14998 17420 15032
rect 17374 14960 17420 14998
rect 17374 14926 17380 14960
rect 17414 14926 17420 14960
rect 17374 14888 17420 14926
rect 17374 14854 17380 14888
rect 17414 14854 17420 14888
rect 17374 14816 17420 14854
rect 17374 14782 17380 14816
rect 17414 14782 17420 14816
rect 17374 14744 17420 14782
rect 17374 14710 17380 14744
rect 17414 14710 17420 14744
rect 17374 14672 17420 14710
rect 17374 14638 17380 14672
rect 17414 14638 17420 14672
rect 17374 14600 17420 14638
rect 17374 14566 17380 14600
rect 17414 14566 17420 14600
rect 17374 14528 17420 14566
rect 17374 14494 17380 14528
rect 17414 14494 17420 14528
rect 17374 14456 17420 14494
rect 17374 14422 17380 14456
rect 17414 14422 17420 14456
rect 17374 14384 17420 14422
rect 17374 14350 17380 14384
rect 17414 14350 17420 14384
rect 17374 14312 17420 14350
rect 17374 14278 17380 14312
rect 17414 14278 17420 14312
rect 17374 14240 17420 14278
rect 17374 14206 17380 14240
rect 17414 14206 17420 14240
rect 17374 14168 17420 14206
rect 17374 14134 17380 14168
rect 17414 14134 17420 14168
rect 17374 14096 17420 14134
rect 17318 14062 17343 14064
rect 17273 14030 17343 14062
rect 17273 13978 17282 14030
rect 17334 13978 17343 14030
rect 17273 13944 17343 13978
rect 17374 14062 17380 14096
rect 17414 14062 17420 14096
rect 17374 14024 17420 14062
rect 17374 13990 17380 14024
rect 17414 13990 17420 14024
rect 17278 13943 17324 13944
rect 17374 13943 17420 13990
rect 17122 13913 17382 13914
rect 13480 13181 13572 13904
rect 16122 13879 16166 13913
rect 16200 13879 16242 13913
rect 13604 13871 13662 13872
rect 13600 13866 13668 13871
rect 13600 13859 13616 13866
rect 13650 13859 13668 13866
rect 13600 13813 13611 13859
rect 13601 13807 13611 13813
rect 13663 13807 13668 13859
rect 14452 13866 15092 13874
rect 14452 13832 14470 13866
rect 14504 13832 14662 13866
rect 14696 13832 14854 13866
rect 14888 13832 15046 13866
rect 15080 13832 15092 13866
rect 14452 13824 15092 13832
rect 13601 13794 13668 13807
rect 16122 13354 16242 13879
rect 17000 13896 17385 13913
rect 17000 13862 17140 13896
rect 17174 13862 17332 13896
rect 17366 13862 17385 13896
rect 17000 13795 17385 13862
rect 16112 13331 16252 13354
rect 16112 13297 16165 13331
rect 16199 13297 16252 13331
rect 16112 13264 16252 13297
rect 17000 13310 17118 13795
rect 17000 13276 17040 13310
rect 17074 13276 17118 13310
rect 17000 13254 17118 13276
rect 13480 13147 13509 13181
rect 13543 13147 13572 13181
rect 13480 13116 13572 13147
rect 13603 13173 13824 13219
rect 13480 13115 13571 13116
rect 13603 13070 13649 13173
rect 13778 13070 13824 13173
rect 13959 13170 14180 13216
rect 13959 13070 14005 13170
rect 14134 13070 14180 13170
rect 14312 13175 14533 13221
rect 14312 13070 14358 13175
rect 14487 13070 14533 13175
rect 14660 13167 14881 13213
rect 13428 13023 13474 13070
rect 13516 13062 13562 13070
rect 13428 12989 13434 13023
rect 13468 12989 13474 13023
rect 13428 12951 13474 12989
rect 13428 12917 13434 12951
rect 13468 12917 13474 12951
rect 13508 13032 13570 13062
rect 13603 13051 13650 13070
rect 13692 13068 13738 13070
rect 13508 12980 13513 13032
rect 13565 12980 13570 13032
rect 13508 12951 13570 12980
rect 13508 12950 13522 12951
rect 13428 12879 13474 12917
rect 13428 12845 13434 12879
rect 13468 12845 13474 12879
rect 13428 12807 13474 12845
rect 13428 12773 13434 12807
rect 13468 12773 13474 12807
rect 13428 12735 13474 12773
rect 13428 12701 13434 12735
rect 13468 12701 13474 12735
rect 13428 12663 13474 12701
rect 13428 12629 13434 12663
rect 13468 12629 13474 12663
rect 13428 12591 13474 12629
rect 13428 12557 13434 12591
rect 13468 12557 13474 12591
rect 13428 12519 13474 12557
rect 13428 12485 13434 12519
rect 13468 12485 13474 12519
rect 13428 12447 13474 12485
rect 13428 12413 13434 12447
rect 13468 12413 13474 12447
rect 13428 12375 13474 12413
rect 13428 12341 13434 12375
rect 13468 12341 13474 12375
rect 13428 12303 13474 12341
rect 13428 12269 13434 12303
rect 13468 12269 13474 12303
rect 13428 12231 13474 12269
rect 13428 12197 13434 12231
rect 13468 12197 13474 12231
rect 13428 12159 13474 12197
rect 13428 12125 13434 12159
rect 13468 12125 13474 12159
rect 13428 12087 13474 12125
rect 13428 12053 13434 12087
rect 13468 12053 13474 12087
rect 13428 12015 13474 12053
rect 13428 11981 13434 12015
rect 13468 11981 13474 12015
rect 13428 11943 13474 11981
rect 13428 11909 13434 11943
rect 13468 11909 13474 11943
rect 13428 11871 13474 11909
rect 13428 11837 13434 11871
rect 13468 11837 13474 11871
rect 13428 11799 13474 11837
rect 13428 11765 13434 11799
rect 13468 11765 13474 11799
rect 13428 11727 13474 11765
rect 13428 11693 13434 11727
rect 13468 11693 13474 11727
rect 13428 11655 13474 11693
rect 13428 11621 13434 11655
rect 13468 11621 13474 11655
rect 13428 11583 13474 11621
rect 13428 11549 13434 11583
rect 13468 11549 13474 11583
rect 13428 11511 13474 11549
rect 13428 11477 13434 11511
rect 13468 11477 13474 11511
rect 13428 11439 13474 11477
rect 13428 11405 13434 11439
rect 13468 11405 13474 11439
rect 13428 11367 13474 11405
rect 13428 11333 13434 11367
rect 13468 11333 13474 11367
rect 13428 11295 13474 11333
rect 13428 11261 13434 11295
rect 13468 11261 13474 11295
rect 13428 11223 13474 11261
rect 13428 11189 13434 11223
rect 13468 11189 13474 11223
rect 13428 11151 13474 11189
rect 13428 11117 13434 11151
rect 13468 11117 13474 11151
rect 13428 10970 13474 11117
rect 13516 12917 13522 12950
rect 13556 12950 13570 12951
rect 13604 13023 13650 13051
rect 13604 12989 13610 13023
rect 13644 12989 13650 13023
rect 13604 12951 13650 12989
rect 13678 13036 13743 13068
rect 13778 13042 13826 13070
rect 13868 13062 13914 13070
rect 13678 12984 13685 13036
rect 13737 12984 13743 13036
rect 13678 12954 13743 12984
rect 13780 13023 13826 13042
rect 13780 12989 13786 13023
rect 13820 12989 13826 13023
rect 13556 12917 13562 12950
rect 13516 12879 13562 12917
rect 13516 12845 13522 12879
rect 13556 12845 13562 12879
rect 13516 12807 13562 12845
rect 13516 12773 13522 12807
rect 13556 12773 13562 12807
rect 13516 12735 13562 12773
rect 13516 12701 13522 12735
rect 13556 12701 13562 12735
rect 13516 12663 13562 12701
rect 13516 12629 13522 12663
rect 13556 12629 13562 12663
rect 13516 12591 13562 12629
rect 13516 12557 13522 12591
rect 13556 12557 13562 12591
rect 13516 12519 13562 12557
rect 13516 12485 13522 12519
rect 13556 12485 13562 12519
rect 13516 12447 13562 12485
rect 13516 12413 13522 12447
rect 13556 12413 13562 12447
rect 13516 12375 13562 12413
rect 13516 12341 13522 12375
rect 13556 12341 13562 12375
rect 13516 12303 13562 12341
rect 13516 12269 13522 12303
rect 13556 12269 13562 12303
rect 13516 12231 13562 12269
rect 13516 12197 13522 12231
rect 13556 12197 13562 12231
rect 13516 12159 13562 12197
rect 13516 12125 13522 12159
rect 13556 12125 13562 12159
rect 13516 12087 13562 12125
rect 13516 12053 13522 12087
rect 13556 12053 13562 12087
rect 13516 12015 13562 12053
rect 13516 11981 13522 12015
rect 13556 11981 13562 12015
rect 13516 11943 13562 11981
rect 13516 11909 13522 11943
rect 13556 11909 13562 11943
rect 13516 11871 13562 11909
rect 13516 11837 13522 11871
rect 13556 11837 13562 11871
rect 13516 11799 13562 11837
rect 13516 11765 13522 11799
rect 13556 11765 13562 11799
rect 13516 11727 13562 11765
rect 13516 11693 13522 11727
rect 13556 11693 13562 11727
rect 13516 11655 13562 11693
rect 13516 11621 13522 11655
rect 13556 11621 13562 11655
rect 13516 11583 13562 11621
rect 13516 11549 13522 11583
rect 13556 11549 13562 11583
rect 13516 11511 13562 11549
rect 13516 11477 13522 11511
rect 13556 11477 13562 11511
rect 13516 11439 13562 11477
rect 13516 11405 13522 11439
rect 13556 11405 13562 11439
rect 13516 11367 13562 11405
rect 13516 11333 13522 11367
rect 13556 11333 13562 11367
rect 13516 11295 13562 11333
rect 13516 11261 13522 11295
rect 13556 11261 13562 11295
rect 13516 11223 13562 11261
rect 13516 11189 13522 11223
rect 13556 11189 13562 11223
rect 13516 11151 13562 11189
rect 13516 11117 13522 11151
rect 13556 11117 13562 11151
rect 13516 11070 13562 11117
rect 13604 12917 13610 12951
rect 13644 12917 13650 12951
rect 13604 12879 13650 12917
rect 13604 12845 13610 12879
rect 13644 12845 13650 12879
rect 13604 12807 13650 12845
rect 13604 12773 13610 12807
rect 13644 12773 13650 12807
rect 13604 12735 13650 12773
rect 13604 12701 13610 12735
rect 13644 12701 13650 12735
rect 13604 12663 13650 12701
rect 13604 12629 13610 12663
rect 13644 12629 13650 12663
rect 13604 12591 13650 12629
rect 13604 12557 13610 12591
rect 13644 12557 13650 12591
rect 13604 12519 13650 12557
rect 13604 12485 13610 12519
rect 13644 12485 13650 12519
rect 13604 12447 13650 12485
rect 13604 12413 13610 12447
rect 13644 12413 13650 12447
rect 13604 12375 13650 12413
rect 13604 12341 13610 12375
rect 13644 12341 13650 12375
rect 13604 12303 13650 12341
rect 13604 12269 13610 12303
rect 13644 12269 13650 12303
rect 13604 12231 13650 12269
rect 13604 12197 13610 12231
rect 13644 12197 13650 12231
rect 13604 12159 13650 12197
rect 13604 12125 13610 12159
rect 13644 12125 13650 12159
rect 13604 12087 13650 12125
rect 13604 12053 13610 12087
rect 13644 12053 13650 12087
rect 13604 12015 13650 12053
rect 13604 11981 13610 12015
rect 13644 11981 13650 12015
rect 13604 11943 13650 11981
rect 13604 11909 13610 11943
rect 13644 11909 13650 11943
rect 13604 11871 13650 11909
rect 13604 11837 13610 11871
rect 13644 11837 13650 11871
rect 13604 11799 13650 11837
rect 13604 11765 13610 11799
rect 13644 11765 13650 11799
rect 13604 11727 13650 11765
rect 13604 11693 13610 11727
rect 13644 11693 13650 11727
rect 13604 11655 13650 11693
rect 13604 11621 13610 11655
rect 13644 11621 13650 11655
rect 13604 11583 13650 11621
rect 13604 11549 13610 11583
rect 13644 11549 13650 11583
rect 13604 11511 13650 11549
rect 13604 11477 13610 11511
rect 13644 11477 13650 11511
rect 13604 11439 13650 11477
rect 13604 11405 13610 11439
rect 13644 11405 13650 11439
rect 13604 11367 13650 11405
rect 13604 11333 13610 11367
rect 13644 11333 13650 11367
rect 13604 11295 13650 11333
rect 13604 11261 13610 11295
rect 13644 11261 13650 11295
rect 13604 11223 13650 11261
rect 13604 11189 13610 11223
rect 13644 11189 13650 11223
rect 13604 11151 13650 11189
rect 13604 11117 13610 11151
rect 13644 11117 13650 11151
rect 13604 11101 13650 11117
rect 13603 11070 13650 11101
rect 13692 12951 13738 12954
rect 13692 12917 13698 12951
rect 13732 12917 13738 12951
rect 13692 12879 13738 12917
rect 13692 12845 13698 12879
rect 13732 12845 13738 12879
rect 13692 12807 13738 12845
rect 13692 12773 13698 12807
rect 13732 12773 13738 12807
rect 13692 12735 13738 12773
rect 13692 12701 13698 12735
rect 13732 12701 13738 12735
rect 13692 12663 13738 12701
rect 13692 12629 13698 12663
rect 13732 12629 13738 12663
rect 13692 12591 13738 12629
rect 13692 12557 13698 12591
rect 13732 12557 13738 12591
rect 13692 12519 13738 12557
rect 13692 12485 13698 12519
rect 13732 12485 13738 12519
rect 13692 12447 13738 12485
rect 13692 12413 13698 12447
rect 13732 12413 13738 12447
rect 13692 12375 13738 12413
rect 13692 12341 13698 12375
rect 13732 12341 13738 12375
rect 13692 12303 13738 12341
rect 13692 12269 13698 12303
rect 13732 12269 13738 12303
rect 13692 12231 13738 12269
rect 13692 12197 13698 12231
rect 13732 12197 13738 12231
rect 13692 12159 13738 12197
rect 13692 12125 13698 12159
rect 13732 12125 13738 12159
rect 13692 12087 13738 12125
rect 13692 12053 13698 12087
rect 13732 12053 13738 12087
rect 13692 12015 13738 12053
rect 13692 11981 13698 12015
rect 13732 11981 13738 12015
rect 13692 11943 13738 11981
rect 13692 11909 13698 11943
rect 13732 11909 13738 11943
rect 13692 11871 13738 11909
rect 13692 11837 13698 11871
rect 13732 11837 13738 11871
rect 13692 11799 13738 11837
rect 13692 11765 13698 11799
rect 13732 11765 13738 11799
rect 13692 11727 13738 11765
rect 13692 11693 13698 11727
rect 13732 11693 13738 11727
rect 13692 11655 13738 11693
rect 13692 11621 13698 11655
rect 13732 11621 13738 11655
rect 13692 11583 13738 11621
rect 13692 11549 13698 11583
rect 13732 11549 13738 11583
rect 13692 11511 13738 11549
rect 13692 11477 13698 11511
rect 13732 11477 13738 11511
rect 13692 11439 13738 11477
rect 13692 11405 13698 11439
rect 13732 11405 13738 11439
rect 13692 11367 13738 11405
rect 13692 11333 13698 11367
rect 13732 11333 13738 11367
rect 13692 11295 13738 11333
rect 13692 11261 13698 11295
rect 13732 11261 13738 11295
rect 13692 11223 13738 11261
rect 13692 11189 13698 11223
rect 13732 11189 13738 11223
rect 13692 11151 13738 11189
rect 13692 11117 13698 11151
rect 13732 11117 13738 11151
rect 13692 11070 13738 11117
rect 13780 12951 13826 12989
rect 13780 12917 13786 12951
rect 13820 12917 13826 12951
rect 13856 13032 13918 13062
rect 13856 12980 13861 13032
rect 13913 12980 13918 13032
rect 13856 12951 13918 12980
rect 13856 12950 13874 12951
rect 13780 12879 13826 12917
rect 13780 12845 13786 12879
rect 13820 12845 13826 12879
rect 13780 12807 13826 12845
rect 13780 12773 13786 12807
rect 13820 12773 13826 12807
rect 13780 12735 13826 12773
rect 13780 12701 13786 12735
rect 13820 12701 13826 12735
rect 13780 12663 13826 12701
rect 13780 12629 13786 12663
rect 13820 12629 13826 12663
rect 13780 12591 13826 12629
rect 13780 12557 13786 12591
rect 13820 12557 13826 12591
rect 13780 12519 13826 12557
rect 13780 12485 13786 12519
rect 13820 12485 13826 12519
rect 13780 12447 13826 12485
rect 13780 12413 13786 12447
rect 13820 12413 13826 12447
rect 13780 12375 13826 12413
rect 13780 12341 13786 12375
rect 13820 12341 13826 12375
rect 13780 12303 13826 12341
rect 13780 12269 13786 12303
rect 13820 12269 13826 12303
rect 13780 12231 13826 12269
rect 13780 12197 13786 12231
rect 13820 12197 13826 12231
rect 13780 12159 13826 12197
rect 13780 12125 13786 12159
rect 13820 12125 13826 12159
rect 13780 12087 13826 12125
rect 13780 12053 13786 12087
rect 13820 12053 13826 12087
rect 13780 12015 13826 12053
rect 13780 11981 13786 12015
rect 13820 11981 13826 12015
rect 13780 11943 13826 11981
rect 13780 11909 13786 11943
rect 13820 11909 13826 11943
rect 13780 11871 13826 11909
rect 13780 11837 13786 11871
rect 13820 11837 13826 11871
rect 13780 11799 13826 11837
rect 13780 11765 13786 11799
rect 13820 11765 13826 11799
rect 13780 11727 13826 11765
rect 13780 11693 13786 11727
rect 13820 11693 13826 11727
rect 13780 11655 13826 11693
rect 13780 11621 13786 11655
rect 13820 11621 13826 11655
rect 13780 11583 13826 11621
rect 13780 11549 13786 11583
rect 13820 11549 13826 11583
rect 13780 11511 13826 11549
rect 13780 11477 13786 11511
rect 13820 11477 13826 11511
rect 13780 11439 13826 11477
rect 13780 11405 13786 11439
rect 13820 11405 13826 11439
rect 13780 11367 13826 11405
rect 13780 11333 13786 11367
rect 13820 11333 13826 11367
rect 13780 11295 13826 11333
rect 13780 11261 13786 11295
rect 13820 11261 13826 11295
rect 13780 11223 13826 11261
rect 13780 11189 13786 11223
rect 13820 11189 13826 11223
rect 13780 11151 13826 11189
rect 13780 11117 13786 11151
rect 13820 11117 13826 11151
rect 13780 11090 13826 11117
rect 13868 12917 13874 12950
rect 13908 12950 13918 12951
rect 13956 13048 14005 13070
rect 13956 13023 14002 13048
rect 13956 12989 13962 13023
rect 13996 12989 14002 13023
rect 13956 12951 14002 12989
rect 14035 13038 14100 13070
rect 14035 12986 14042 13038
rect 14094 12986 14100 13038
rect 14035 12956 14100 12986
rect 14132 13039 14180 13070
rect 14220 13068 14266 13070
rect 14132 13023 14178 13039
rect 14132 12989 14138 13023
rect 14172 12989 14178 13023
rect 13908 12917 13914 12950
rect 13868 12879 13914 12917
rect 13868 12845 13874 12879
rect 13908 12845 13914 12879
rect 13868 12807 13914 12845
rect 13868 12773 13874 12807
rect 13908 12773 13914 12807
rect 13868 12735 13914 12773
rect 13868 12701 13874 12735
rect 13908 12701 13914 12735
rect 13868 12663 13914 12701
rect 13868 12629 13874 12663
rect 13908 12629 13914 12663
rect 13868 12591 13914 12629
rect 13868 12557 13874 12591
rect 13908 12557 13914 12591
rect 13868 12519 13914 12557
rect 13868 12485 13874 12519
rect 13908 12485 13914 12519
rect 13868 12447 13914 12485
rect 13868 12413 13874 12447
rect 13908 12413 13914 12447
rect 13868 12375 13914 12413
rect 13868 12341 13874 12375
rect 13908 12341 13914 12375
rect 13868 12303 13914 12341
rect 13868 12269 13874 12303
rect 13908 12269 13914 12303
rect 13868 12231 13914 12269
rect 13868 12197 13874 12231
rect 13908 12197 13914 12231
rect 13868 12159 13914 12197
rect 13868 12125 13874 12159
rect 13908 12125 13914 12159
rect 13868 12087 13914 12125
rect 13868 12053 13874 12087
rect 13908 12053 13914 12087
rect 13868 12015 13914 12053
rect 13868 11981 13874 12015
rect 13908 11981 13914 12015
rect 13868 11943 13914 11981
rect 13868 11909 13874 11943
rect 13908 11909 13914 11943
rect 13868 11871 13914 11909
rect 13868 11837 13874 11871
rect 13908 11837 13914 11871
rect 13868 11799 13914 11837
rect 13868 11765 13874 11799
rect 13908 11765 13914 11799
rect 13868 11727 13914 11765
rect 13868 11693 13874 11727
rect 13908 11693 13914 11727
rect 13868 11655 13914 11693
rect 13868 11621 13874 11655
rect 13908 11621 13914 11655
rect 13868 11583 13914 11621
rect 13868 11549 13874 11583
rect 13908 11549 13914 11583
rect 13868 11511 13914 11549
rect 13868 11477 13874 11511
rect 13908 11477 13914 11511
rect 13868 11439 13914 11477
rect 13868 11405 13874 11439
rect 13908 11405 13914 11439
rect 13868 11367 13914 11405
rect 13868 11333 13874 11367
rect 13908 11333 13914 11367
rect 13868 11295 13914 11333
rect 13868 11261 13874 11295
rect 13908 11261 13914 11295
rect 13868 11223 13914 11261
rect 13868 11189 13874 11223
rect 13908 11189 13914 11223
rect 13868 11151 13914 11189
rect 13868 11117 13874 11151
rect 13908 11117 13914 11151
rect 13780 11070 13827 11090
rect 13868 11070 13914 11117
rect 13956 12917 13962 12951
rect 13996 12917 14002 12951
rect 13956 12879 14002 12917
rect 13956 12845 13962 12879
rect 13996 12845 14002 12879
rect 13956 12807 14002 12845
rect 13956 12773 13962 12807
rect 13996 12773 14002 12807
rect 13956 12735 14002 12773
rect 13956 12701 13962 12735
rect 13996 12701 14002 12735
rect 13956 12663 14002 12701
rect 13956 12629 13962 12663
rect 13996 12629 14002 12663
rect 13956 12591 14002 12629
rect 13956 12557 13962 12591
rect 13996 12557 14002 12591
rect 13956 12519 14002 12557
rect 13956 12485 13962 12519
rect 13996 12485 14002 12519
rect 13956 12447 14002 12485
rect 13956 12413 13962 12447
rect 13996 12413 14002 12447
rect 13956 12375 14002 12413
rect 13956 12341 13962 12375
rect 13996 12341 14002 12375
rect 13956 12303 14002 12341
rect 13956 12269 13962 12303
rect 13996 12269 14002 12303
rect 13956 12231 14002 12269
rect 13956 12197 13962 12231
rect 13996 12197 14002 12231
rect 13956 12159 14002 12197
rect 13956 12125 13962 12159
rect 13996 12125 14002 12159
rect 13956 12087 14002 12125
rect 13956 12053 13962 12087
rect 13996 12053 14002 12087
rect 13956 12015 14002 12053
rect 13956 11981 13962 12015
rect 13996 11981 14002 12015
rect 13956 11943 14002 11981
rect 13956 11909 13962 11943
rect 13996 11909 14002 11943
rect 13956 11871 14002 11909
rect 13956 11837 13962 11871
rect 13996 11837 14002 11871
rect 13956 11799 14002 11837
rect 13956 11765 13962 11799
rect 13996 11765 14002 11799
rect 13956 11727 14002 11765
rect 13956 11693 13962 11727
rect 13996 11693 14002 11727
rect 13956 11655 14002 11693
rect 13956 11621 13962 11655
rect 13996 11621 14002 11655
rect 13956 11583 14002 11621
rect 13956 11549 13962 11583
rect 13996 11549 14002 11583
rect 13956 11511 14002 11549
rect 13956 11477 13962 11511
rect 13996 11477 14002 11511
rect 13956 11439 14002 11477
rect 13956 11405 13962 11439
rect 13996 11405 14002 11439
rect 13956 11367 14002 11405
rect 13956 11333 13962 11367
rect 13996 11333 14002 11367
rect 13956 11295 14002 11333
rect 13956 11261 13962 11295
rect 13996 11261 14002 11295
rect 13956 11223 14002 11261
rect 13956 11189 13962 11223
rect 13996 11189 14002 11223
rect 13956 11151 14002 11189
rect 13956 11117 13962 11151
rect 13996 11117 14002 11151
rect 13603 10970 13649 11070
rect 13428 10924 13649 10970
rect 13781 10968 13827 11070
rect 13956 10968 14002 11117
rect 14044 12951 14090 12956
rect 14044 12917 14050 12951
rect 14084 12917 14090 12951
rect 14044 12879 14090 12917
rect 14044 12845 14050 12879
rect 14084 12845 14090 12879
rect 14044 12807 14090 12845
rect 14044 12773 14050 12807
rect 14084 12773 14090 12807
rect 14044 12735 14090 12773
rect 14044 12701 14050 12735
rect 14084 12701 14090 12735
rect 14044 12663 14090 12701
rect 14044 12629 14050 12663
rect 14084 12629 14090 12663
rect 14044 12591 14090 12629
rect 14044 12557 14050 12591
rect 14084 12557 14090 12591
rect 14044 12519 14090 12557
rect 14044 12485 14050 12519
rect 14084 12485 14090 12519
rect 14044 12447 14090 12485
rect 14044 12413 14050 12447
rect 14084 12413 14090 12447
rect 14044 12375 14090 12413
rect 14044 12341 14050 12375
rect 14084 12341 14090 12375
rect 14044 12303 14090 12341
rect 14044 12269 14050 12303
rect 14084 12269 14090 12303
rect 14044 12231 14090 12269
rect 14044 12197 14050 12231
rect 14084 12197 14090 12231
rect 14044 12159 14090 12197
rect 14044 12125 14050 12159
rect 14084 12125 14090 12159
rect 14044 12087 14090 12125
rect 14044 12053 14050 12087
rect 14084 12053 14090 12087
rect 14044 12015 14090 12053
rect 14044 11981 14050 12015
rect 14084 11981 14090 12015
rect 14044 11943 14090 11981
rect 14044 11909 14050 11943
rect 14084 11909 14090 11943
rect 14044 11871 14090 11909
rect 14044 11837 14050 11871
rect 14084 11837 14090 11871
rect 14044 11799 14090 11837
rect 14044 11765 14050 11799
rect 14084 11765 14090 11799
rect 14044 11727 14090 11765
rect 14044 11693 14050 11727
rect 14084 11693 14090 11727
rect 14044 11655 14090 11693
rect 14044 11621 14050 11655
rect 14084 11621 14090 11655
rect 14044 11583 14090 11621
rect 14044 11549 14050 11583
rect 14084 11549 14090 11583
rect 14044 11511 14090 11549
rect 14044 11477 14050 11511
rect 14084 11477 14090 11511
rect 14044 11439 14090 11477
rect 14044 11405 14050 11439
rect 14084 11405 14090 11439
rect 14044 11367 14090 11405
rect 14044 11333 14050 11367
rect 14084 11333 14090 11367
rect 14044 11295 14090 11333
rect 14044 11261 14050 11295
rect 14084 11261 14090 11295
rect 14044 11223 14090 11261
rect 14044 11189 14050 11223
rect 14084 11189 14090 11223
rect 14044 11151 14090 11189
rect 14044 11117 14050 11151
rect 14084 11117 14090 11151
rect 14044 11070 14090 11117
rect 14132 12951 14178 12989
rect 14212 13038 14274 13068
rect 14212 12986 14217 13038
rect 14269 12986 14274 13038
rect 14212 12956 14274 12986
rect 14308 13053 14358 13070
rect 14308 13023 14354 13053
rect 14308 12989 14314 13023
rect 14348 12989 14354 13023
rect 14132 12917 14138 12951
rect 14172 12917 14178 12951
rect 14132 12879 14178 12917
rect 14132 12845 14138 12879
rect 14172 12845 14178 12879
rect 14132 12807 14178 12845
rect 14132 12773 14138 12807
rect 14172 12773 14178 12807
rect 14132 12735 14178 12773
rect 14132 12701 14138 12735
rect 14172 12701 14178 12735
rect 14132 12663 14178 12701
rect 14132 12629 14138 12663
rect 14172 12629 14178 12663
rect 14132 12591 14178 12629
rect 14132 12557 14138 12591
rect 14172 12557 14178 12591
rect 14132 12519 14178 12557
rect 14132 12485 14138 12519
rect 14172 12485 14178 12519
rect 14132 12447 14178 12485
rect 14132 12413 14138 12447
rect 14172 12413 14178 12447
rect 14132 12375 14178 12413
rect 14132 12341 14138 12375
rect 14172 12341 14178 12375
rect 14132 12303 14178 12341
rect 14132 12269 14138 12303
rect 14172 12269 14178 12303
rect 14132 12231 14178 12269
rect 14132 12197 14138 12231
rect 14172 12197 14178 12231
rect 14132 12159 14178 12197
rect 14132 12125 14138 12159
rect 14172 12125 14178 12159
rect 14132 12087 14178 12125
rect 14132 12053 14138 12087
rect 14172 12053 14178 12087
rect 14132 12015 14178 12053
rect 14132 11981 14138 12015
rect 14172 11981 14178 12015
rect 14132 11943 14178 11981
rect 14132 11909 14138 11943
rect 14172 11909 14178 11943
rect 14132 11871 14178 11909
rect 14132 11837 14138 11871
rect 14172 11837 14178 11871
rect 14132 11799 14178 11837
rect 14132 11765 14138 11799
rect 14172 11765 14178 11799
rect 14132 11727 14178 11765
rect 14132 11693 14138 11727
rect 14172 11693 14178 11727
rect 14132 11655 14178 11693
rect 14132 11621 14138 11655
rect 14172 11621 14178 11655
rect 14132 11583 14178 11621
rect 14132 11549 14138 11583
rect 14172 11549 14178 11583
rect 14132 11511 14178 11549
rect 14132 11477 14138 11511
rect 14172 11477 14178 11511
rect 14132 11439 14178 11477
rect 14132 11405 14138 11439
rect 14172 11405 14178 11439
rect 14132 11367 14178 11405
rect 14132 11333 14138 11367
rect 14172 11333 14178 11367
rect 14132 11295 14178 11333
rect 14132 11261 14138 11295
rect 14172 11261 14178 11295
rect 14132 11223 14178 11261
rect 14132 11189 14138 11223
rect 14172 11189 14178 11223
rect 14132 11151 14178 11189
rect 14132 11117 14138 11151
rect 14172 11117 14178 11151
rect 13781 10922 14002 10968
rect 14132 10970 14178 11117
rect 14220 12951 14266 12956
rect 14220 12917 14226 12951
rect 14260 12917 14266 12951
rect 14220 12879 14266 12917
rect 14220 12845 14226 12879
rect 14260 12845 14266 12879
rect 14220 12807 14266 12845
rect 14220 12773 14226 12807
rect 14260 12773 14266 12807
rect 14220 12735 14266 12773
rect 14220 12701 14226 12735
rect 14260 12701 14266 12735
rect 14220 12663 14266 12701
rect 14220 12629 14226 12663
rect 14260 12629 14266 12663
rect 14220 12591 14266 12629
rect 14220 12557 14226 12591
rect 14260 12557 14266 12591
rect 14220 12519 14266 12557
rect 14220 12485 14226 12519
rect 14260 12485 14266 12519
rect 14220 12447 14266 12485
rect 14220 12413 14226 12447
rect 14260 12413 14266 12447
rect 14220 12375 14266 12413
rect 14220 12341 14226 12375
rect 14260 12341 14266 12375
rect 14220 12303 14266 12341
rect 14220 12269 14226 12303
rect 14260 12269 14266 12303
rect 14220 12231 14266 12269
rect 14220 12197 14226 12231
rect 14260 12197 14266 12231
rect 14220 12159 14266 12197
rect 14220 12125 14226 12159
rect 14260 12125 14266 12159
rect 14220 12087 14266 12125
rect 14220 12053 14226 12087
rect 14260 12053 14266 12087
rect 14220 12015 14266 12053
rect 14220 11981 14226 12015
rect 14260 11981 14266 12015
rect 14220 11943 14266 11981
rect 14220 11909 14226 11943
rect 14260 11909 14266 11943
rect 14220 11871 14266 11909
rect 14220 11837 14226 11871
rect 14260 11837 14266 11871
rect 14220 11799 14266 11837
rect 14220 11765 14226 11799
rect 14260 11765 14266 11799
rect 14220 11727 14266 11765
rect 14220 11693 14226 11727
rect 14260 11693 14266 11727
rect 14220 11655 14266 11693
rect 14220 11621 14226 11655
rect 14260 11621 14266 11655
rect 14220 11583 14266 11621
rect 14220 11549 14226 11583
rect 14260 11549 14266 11583
rect 14220 11511 14266 11549
rect 14220 11477 14226 11511
rect 14260 11477 14266 11511
rect 14220 11439 14266 11477
rect 14220 11405 14226 11439
rect 14260 11405 14266 11439
rect 14220 11367 14266 11405
rect 14220 11333 14226 11367
rect 14260 11333 14266 11367
rect 14220 11295 14266 11333
rect 14220 11261 14226 11295
rect 14260 11261 14266 11295
rect 14220 11223 14266 11261
rect 14220 11189 14226 11223
rect 14260 11189 14266 11223
rect 14220 11151 14266 11189
rect 14220 11117 14226 11151
rect 14260 11117 14266 11151
rect 14220 11070 14266 11117
rect 14308 12951 14354 12989
rect 14388 13038 14453 13070
rect 14388 12986 14395 13038
rect 14447 12986 14453 13038
rect 14388 12956 14453 12986
rect 14484 13044 14533 13070
rect 14572 13066 14618 13070
rect 14484 13023 14530 13044
rect 14484 12989 14490 13023
rect 14524 12989 14530 13023
rect 14308 12917 14314 12951
rect 14348 12917 14354 12951
rect 14308 12879 14354 12917
rect 14308 12845 14314 12879
rect 14348 12845 14354 12879
rect 14308 12807 14354 12845
rect 14308 12773 14314 12807
rect 14348 12773 14354 12807
rect 14308 12735 14354 12773
rect 14308 12701 14314 12735
rect 14348 12701 14354 12735
rect 14308 12663 14354 12701
rect 14308 12629 14314 12663
rect 14348 12629 14354 12663
rect 14308 12591 14354 12629
rect 14308 12557 14314 12591
rect 14348 12557 14354 12591
rect 14308 12519 14354 12557
rect 14308 12485 14314 12519
rect 14348 12485 14354 12519
rect 14308 12447 14354 12485
rect 14308 12413 14314 12447
rect 14348 12413 14354 12447
rect 14308 12375 14354 12413
rect 14308 12341 14314 12375
rect 14348 12341 14354 12375
rect 14308 12303 14354 12341
rect 14308 12269 14314 12303
rect 14348 12269 14354 12303
rect 14308 12231 14354 12269
rect 14308 12197 14314 12231
rect 14348 12197 14354 12231
rect 14308 12159 14354 12197
rect 14308 12125 14314 12159
rect 14348 12125 14354 12159
rect 14308 12087 14354 12125
rect 14308 12053 14314 12087
rect 14348 12053 14354 12087
rect 14308 12015 14354 12053
rect 14308 11981 14314 12015
rect 14348 11981 14354 12015
rect 14308 11943 14354 11981
rect 14308 11909 14314 11943
rect 14348 11909 14354 11943
rect 14308 11871 14354 11909
rect 14308 11837 14314 11871
rect 14348 11837 14354 11871
rect 14308 11799 14354 11837
rect 14308 11765 14314 11799
rect 14348 11765 14354 11799
rect 14308 11727 14354 11765
rect 14308 11693 14314 11727
rect 14348 11693 14354 11727
rect 14308 11655 14354 11693
rect 14308 11621 14314 11655
rect 14348 11621 14354 11655
rect 14308 11583 14354 11621
rect 14308 11549 14314 11583
rect 14348 11549 14354 11583
rect 14308 11511 14354 11549
rect 14308 11477 14314 11511
rect 14348 11477 14354 11511
rect 14308 11439 14354 11477
rect 14308 11405 14314 11439
rect 14348 11405 14354 11439
rect 14308 11367 14354 11405
rect 14308 11333 14314 11367
rect 14348 11333 14354 11367
rect 14308 11295 14354 11333
rect 14308 11261 14314 11295
rect 14348 11261 14354 11295
rect 14308 11223 14354 11261
rect 14308 11189 14314 11223
rect 14348 11189 14354 11223
rect 14308 11151 14354 11189
rect 14308 11117 14314 11151
rect 14348 11117 14354 11151
rect 14308 11101 14354 11117
rect 14307 11070 14354 11101
rect 14396 12951 14442 12956
rect 14396 12917 14402 12951
rect 14436 12917 14442 12951
rect 14396 12879 14442 12917
rect 14396 12845 14402 12879
rect 14436 12845 14442 12879
rect 14396 12807 14442 12845
rect 14396 12773 14402 12807
rect 14436 12773 14442 12807
rect 14396 12735 14442 12773
rect 14396 12701 14402 12735
rect 14436 12701 14442 12735
rect 14396 12663 14442 12701
rect 14396 12629 14402 12663
rect 14436 12629 14442 12663
rect 14396 12591 14442 12629
rect 14396 12557 14402 12591
rect 14436 12557 14442 12591
rect 14396 12519 14442 12557
rect 14396 12485 14402 12519
rect 14436 12485 14442 12519
rect 14396 12447 14442 12485
rect 14396 12413 14402 12447
rect 14436 12413 14442 12447
rect 14396 12375 14442 12413
rect 14396 12341 14402 12375
rect 14436 12341 14442 12375
rect 14396 12303 14442 12341
rect 14396 12269 14402 12303
rect 14436 12269 14442 12303
rect 14396 12231 14442 12269
rect 14396 12197 14402 12231
rect 14436 12197 14442 12231
rect 14396 12159 14442 12197
rect 14396 12125 14402 12159
rect 14436 12125 14442 12159
rect 14396 12087 14442 12125
rect 14396 12053 14402 12087
rect 14436 12053 14442 12087
rect 14396 12015 14442 12053
rect 14396 11981 14402 12015
rect 14436 11981 14442 12015
rect 14396 11943 14442 11981
rect 14396 11909 14402 11943
rect 14436 11909 14442 11943
rect 14396 11871 14442 11909
rect 14396 11837 14402 11871
rect 14436 11837 14442 11871
rect 14396 11799 14442 11837
rect 14396 11765 14402 11799
rect 14436 11765 14442 11799
rect 14396 11727 14442 11765
rect 14396 11693 14402 11727
rect 14436 11693 14442 11727
rect 14396 11655 14442 11693
rect 14396 11621 14402 11655
rect 14436 11621 14442 11655
rect 14396 11583 14442 11621
rect 14396 11549 14402 11583
rect 14436 11549 14442 11583
rect 14396 11511 14442 11549
rect 14396 11477 14402 11511
rect 14436 11477 14442 11511
rect 14396 11439 14442 11477
rect 14396 11405 14402 11439
rect 14436 11405 14442 11439
rect 14396 11367 14442 11405
rect 14396 11333 14402 11367
rect 14436 11333 14442 11367
rect 14396 11295 14442 11333
rect 14396 11261 14402 11295
rect 14436 11261 14442 11295
rect 14396 11223 14442 11261
rect 14396 11189 14402 11223
rect 14436 11189 14442 11223
rect 14396 11151 14442 11189
rect 14396 11117 14402 11151
rect 14436 11117 14442 11151
rect 14396 11070 14442 11117
rect 14484 12951 14530 12989
rect 14562 13036 14624 13066
rect 14562 12984 14567 13036
rect 14619 12984 14624 13036
rect 14562 12954 14624 12984
rect 14660 13023 14706 13167
rect 14660 12989 14666 13023
rect 14700 12989 14706 13023
rect 14484 12917 14490 12951
rect 14524 12917 14530 12951
rect 14484 12879 14530 12917
rect 14484 12845 14490 12879
rect 14524 12845 14530 12879
rect 14484 12807 14530 12845
rect 14484 12773 14490 12807
rect 14524 12773 14530 12807
rect 14484 12735 14530 12773
rect 14484 12701 14490 12735
rect 14524 12701 14530 12735
rect 14484 12663 14530 12701
rect 14484 12629 14490 12663
rect 14524 12629 14530 12663
rect 14484 12591 14530 12629
rect 14484 12557 14490 12591
rect 14524 12557 14530 12591
rect 14484 12519 14530 12557
rect 14484 12485 14490 12519
rect 14524 12485 14530 12519
rect 14484 12447 14530 12485
rect 14484 12413 14490 12447
rect 14524 12413 14530 12447
rect 14484 12375 14530 12413
rect 14484 12341 14490 12375
rect 14524 12341 14530 12375
rect 14484 12303 14530 12341
rect 14484 12269 14490 12303
rect 14524 12269 14530 12303
rect 14484 12231 14530 12269
rect 14484 12197 14490 12231
rect 14524 12197 14530 12231
rect 14484 12159 14530 12197
rect 14484 12125 14490 12159
rect 14524 12125 14530 12159
rect 14484 12087 14530 12125
rect 14484 12053 14490 12087
rect 14524 12053 14530 12087
rect 14484 12015 14530 12053
rect 14484 11981 14490 12015
rect 14524 11981 14530 12015
rect 14484 11943 14530 11981
rect 14484 11909 14490 11943
rect 14524 11909 14530 11943
rect 14484 11871 14530 11909
rect 14484 11837 14490 11871
rect 14524 11837 14530 11871
rect 14484 11799 14530 11837
rect 14484 11765 14490 11799
rect 14524 11765 14530 11799
rect 14484 11727 14530 11765
rect 14484 11693 14490 11727
rect 14524 11693 14530 11727
rect 14484 11655 14530 11693
rect 14484 11621 14490 11655
rect 14524 11621 14530 11655
rect 14484 11583 14530 11621
rect 14484 11549 14490 11583
rect 14524 11549 14530 11583
rect 14484 11511 14530 11549
rect 14484 11477 14490 11511
rect 14524 11477 14530 11511
rect 14484 11439 14530 11477
rect 14484 11405 14490 11439
rect 14524 11405 14530 11439
rect 14484 11367 14530 11405
rect 14484 11333 14490 11367
rect 14524 11333 14530 11367
rect 14484 11295 14530 11333
rect 14484 11261 14490 11295
rect 14524 11261 14530 11295
rect 14484 11223 14530 11261
rect 14484 11189 14490 11223
rect 14524 11189 14530 11223
rect 14484 11151 14530 11189
rect 14484 11117 14490 11151
rect 14524 11117 14530 11151
rect 14307 10970 14353 11070
rect 14484 10994 14530 11117
rect 14572 12951 14618 12954
rect 14572 12917 14578 12951
rect 14612 12917 14618 12951
rect 14572 12879 14618 12917
rect 14572 12845 14578 12879
rect 14612 12845 14618 12879
rect 14572 12807 14618 12845
rect 14572 12773 14578 12807
rect 14612 12773 14618 12807
rect 14572 12735 14618 12773
rect 14572 12701 14578 12735
rect 14612 12701 14618 12735
rect 14572 12663 14618 12701
rect 14572 12629 14578 12663
rect 14612 12629 14618 12663
rect 14572 12591 14618 12629
rect 14572 12557 14578 12591
rect 14612 12557 14618 12591
rect 14572 12519 14618 12557
rect 14572 12485 14578 12519
rect 14612 12485 14618 12519
rect 14572 12447 14618 12485
rect 14572 12413 14578 12447
rect 14612 12413 14618 12447
rect 14572 12375 14618 12413
rect 14572 12341 14578 12375
rect 14612 12341 14618 12375
rect 14572 12303 14618 12341
rect 14572 12269 14578 12303
rect 14612 12269 14618 12303
rect 14572 12231 14618 12269
rect 14572 12197 14578 12231
rect 14612 12197 14618 12231
rect 14572 12159 14618 12197
rect 14572 12125 14578 12159
rect 14612 12125 14618 12159
rect 14572 12087 14618 12125
rect 14572 12053 14578 12087
rect 14612 12053 14618 12087
rect 14572 12015 14618 12053
rect 14572 11981 14578 12015
rect 14612 11981 14618 12015
rect 14572 11943 14618 11981
rect 14572 11909 14578 11943
rect 14612 11909 14618 11943
rect 14572 11871 14618 11909
rect 14572 11837 14578 11871
rect 14612 11837 14618 11871
rect 14572 11799 14618 11837
rect 14572 11765 14578 11799
rect 14612 11765 14618 11799
rect 14572 11727 14618 11765
rect 14572 11693 14578 11727
rect 14612 11693 14618 11727
rect 14572 11655 14618 11693
rect 14572 11621 14578 11655
rect 14612 11621 14618 11655
rect 14572 11583 14618 11621
rect 14572 11549 14578 11583
rect 14612 11549 14618 11583
rect 14572 11511 14618 11549
rect 14572 11477 14578 11511
rect 14612 11477 14618 11511
rect 14572 11439 14618 11477
rect 14572 11405 14578 11439
rect 14612 11405 14618 11439
rect 14572 11367 14618 11405
rect 14572 11333 14578 11367
rect 14612 11333 14618 11367
rect 14572 11295 14618 11333
rect 14572 11261 14578 11295
rect 14612 11261 14618 11295
rect 14572 11223 14618 11261
rect 14572 11189 14578 11223
rect 14612 11189 14618 11223
rect 14572 11151 14618 11189
rect 14572 11117 14578 11151
rect 14612 11117 14618 11151
rect 14572 11070 14618 11117
rect 14660 12951 14706 12989
rect 14740 13039 14805 13071
rect 14740 12987 14747 13039
rect 14799 12987 14805 13039
rect 14835 13070 14881 13167
rect 15016 13175 15237 13221
rect 15016 13070 15062 13175
rect 15191 13070 15237 13175
rect 15366 13175 15587 13221
rect 15366 13070 15412 13175
rect 15541 13070 15587 13175
rect 15720 13173 15941 13219
rect 15720 13070 15766 13173
rect 15895 13070 15941 13173
rect 16069 13171 16290 13217
rect 16069 13070 16115 13171
rect 14835 13036 14882 13070
rect 14924 13066 14970 13070
rect 14740 12957 14805 12987
rect 14836 13023 14882 13036
rect 14836 12989 14842 13023
rect 14876 12989 14882 13023
rect 14660 12917 14666 12951
rect 14700 12917 14706 12951
rect 14660 12879 14706 12917
rect 14660 12845 14666 12879
rect 14700 12845 14706 12879
rect 14660 12807 14706 12845
rect 14660 12773 14666 12807
rect 14700 12773 14706 12807
rect 14660 12735 14706 12773
rect 14660 12701 14666 12735
rect 14700 12701 14706 12735
rect 14660 12663 14706 12701
rect 14660 12629 14666 12663
rect 14700 12629 14706 12663
rect 14660 12591 14706 12629
rect 14660 12557 14666 12591
rect 14700 12557 14706 12591
rect 14660 12519 14706 12557
rect 14660 12485 14666 12519
rect 14700 12485 14706 12519
rect 14660 12447 14706 12485
rect 14660 12413 14666 12447
rect 14700 12413 14706 12447
rect 14660 12375 14706 12413
rect 14660 12341 14666 12375
rect 14700 12341 14706 12375
rect 14660 12303 14706 12341
rect 14660 12269 14666 12303
rect 14700 12269 14706 12303
rect 14660 12231 14706 12269
rect 14660 12197 14666 12231
rect 14700 12197 14706 12231
rect 14660 12159 14706 12197
rect 14660 12125 14666 12159
rect 14700 12125 14706 12159
rect 14660 12087 14706 12125
rect 14660 12053 14666 12087
rect 14700 12053 14706 12087
rect 14660 12015 14706 12053
rect 14660 11981 14666 12015
rect 14700 11981 14706 12015
rect 14660 11943 14706 11981
rect 14660 11909 14666 11943
rect 14700 11909 14706 11943
rect 14660 11871 14706 11909
rect 14660 11837 14666 11871
rect 14700 11837 14706 11871
rect 14660 11799 14706 11837
rect 14660 11765 14666 11799
rect 14700 11765 14706 11799
rect 14660 11727 14706 11765
rect 14660 11693 14666 11727
rect 14700 11693 14706 11727
rect 14660 11655 14706 11693
rect 14660 11621 14666 11655
rect 14700 11621 14706 11655
rect 14660 11583 14706 11621
rect 14660 11549 14666 11583
rect 14700 11549 14706 11583
rect 14660 11511 14706 11549
rect 14660 11477 14666 11511
rect 14700 11477 14706 11511
rect 14660 11439 14706 11477
rect 14660 11405 14666 11439
rect 14700 11405 14706 11439
rect 14660 11367 14706 11405
rect 14660 11333 14666 11367
rect 14700 11333 14706 11367
rect 14660 11295 14706 11333
rect 14660 11261 14666 11295
rect 14700 11261 14706 11295
rect 14660 11223 14706 11261
rect 14660 11189 14666 11223
rect 14700 11189 14706 11223
rect 14660 11151 14706 11189
rect 14660 11117 14666 11151
rect 14700 11117 14706 11151
rect 14660 11101 14706 11117
rect 14659 11070 14706 11101
rect 14748 12951 14794 12957
rect 14748 12917 14754 12951
rect 14788 12917 14794 12951
rect 14748 12879 14794 12917
rect 14748 12845 14754 12879
rect 14788 12845 14794 12879
rect 14748 12807 14794 12845
rect 14748 12773 14754 12807
rect 14788 12773 14794 12807
rect 14748 12735 14794 12773
rect 14748 12701 14754 12735
rect 14788 12701 14794 12735
rect 14748 12663 14794 12701
rect 14748 12629 14754 12663
rect 14788 12629 14794 12663
rect 14748 12591 14794 12629
rect 14748 12557 14754 12591
rect 14788 12557 14794 12591
rect 14748 12519 14794 12557
rect 14748 12485 14754 12519
rect 14788 12485 14794 12519
rect 14748 12447 14794 12485
rect 14748 12413 14754 12447
rect 14788 12413 14794 12447
rect 14748 12375 14794 12413
rect 14748 12341 14754 12375
rect 14788 12341 14794 12375
rect 14748 12303 14794 12341
rect 14748 12269 14754 12303
rect 14788 12269 14794 12303
rect 14748 12231 14794 12269
rect 14748 12197 14754 12231
rect 14788 12197 14794 12231
rect 14748 12159 14794 12197
rect 14748 12125 14754 12159
rect 14788 12125 14794 12159
rect 14748 12087 14794 12125
rect 14748 12053 14754 12087
rect 14788 12053 14794 12087
rect 14748 12015 14794 12053
rect 14748 11981 14754 12015
rect 14788 11981 14794 12015
rect 14748 11943 14794 11981
rect 14748 11909 14754 11943
rect 14788 11909 14794 11943
rect 14748 11871 14794 11909
rect 14748 11837 14754 11871
rect 14788 11837 14794 11871
rect 14748 11799 14794 11837
rect 14748 11765 14754 11799
rect 14788 11765 14794 11799
rect 14748 11727 14794 11765
rect 14748 11693 14754 11727
rect 14788 11693 14794 11727
rect 14748 11655 14794 11693
rect 14748 11621 14754 11655
rect 14788 11621 14794 11655
rect 14748 11583 14794 11621
rect 14748 11549 14754 11583
rect 14788 11549 14794 11583
rect 14748 11511 14794 11549
rect 14748 11477 14754 11511
rect 14788 11477 14794 11511
rect 14748 11439 14794 11477
rect 14748 11405 14754 11439
rect 14788 11405 14794 11439
rect 14748 11367 14794 11405
rect 14748 11333 14754 11367
rect 14788 11333 14794 11367
rect 14748 11295 14794 11333
rect 14748 11261 14754 11295
rect 14788 11261 14794 11295
rect 14748 11223 14794 11261
rect 14748 11189 14754 11223
rect 14788 11189 14794 11223
rect 14748 11151 14794 11189
rect 14748 11117 14754 11151
rect 14788 11117 14794 11151
rect 14748 11070 14794 11117
rect 14836 12951 14882 12989
rect 14916 13036 14978 13066
rect 14916 12984 14921 13036
rect 14973 12984 14978 13036
rect 14916 12954 14978 12984
rect 15012 13053 15062 13070
rect 15012 13023 15058 13053
rect 15012 12989 15018 13023
rect 15052 12989 15058 13023
rect 14836 12917 14842 12951
rect 14876 12917 14882 12951
rect 14836 12879 14882 12917
rect 14836 12845 14842 12879
rect 14876 12845 14882 12879
rect 14836 12807 14882 12845
rect 14836 12773 14842 12807
rect 14876 12773 14882 12807
rect 14836 12735 14882 12773
rect 14836 12701 14842 12735
rect 14876 12701 14882 12735
rect 14836 12663 14882 12701
rect 14836 12629 14842 12663
rect 14876 12629 14882 12663
rect 14836 12591 14882 12629
rect 14836 12557 14842 12591
rect 14876 12557 14882 12591
rect 14836 12519 14882 12557
rect 14836 12485 14842 12519
rect 14876 12485 14882 12519
rect 14836 12447 14882 12485
rect 14836 12413 14842 12447
rect 14876 12413 14882 12447
rect 14836 12375 14882 12413
rect 14836 12341 14842 12375
rect 14876 12341 14882 12375
rect 14836 12303 14882 12341
rect 14836 12269 14842 12303
rect 14876 12269 14882 12303
rect 14836 12231 14882 12269
rect 14836 12197 14842 12231
rect 14876 12197 14882 12231
rect 14836 12159 14882 12197
rect 14836 12125 14842 12159
rect 14876 12125 14882 12159
rect 14836 12087 14882 12125
rect 14836 12053 14842 12087
rect 14876 12053 14882 12087
rect 14836 12015 14882 12053
rect 14836 11981 14842 12015
rect 14876 11981 14882 12015
rect 14836 11943 14882 11981
rect 14836 11909 14842 11943
rect 14876 11909 14882 11943
rect 14836 11871 14882 11909
rect 14836 11837 14842 11871
rect 14876 11837 14882 11871
rect 14836 11799 14882 11837
rect 14836 11765 14842 11799
rect 14876 11765 14882 11799
rect 14836 11727 14882 11765
rect 14836 11693 14842 11727
rect 14876 11693 14882 11727
rect 14836 11655 14882 11693
rect 14836 11621 14842 11655
rect 14876 11621 14882 11655
rect 14836 11583 14882 11621
rect 14836 11549 14842 11583
rect 14876 11549 14882 11583
rect 14836 11511 14882 11549
rect 14836 11477 14842 11511
rect 14876 11477 14882 11511
rect 14836 11439 14882 11477
rect 14836 11405 14842 11439
rect 14876 11405 14882 11439
rect 14836 11367 14882 11405
rect 14836 11333 14842 11367
rect 14876 11333 14882 11367
rect 14836 11295 14882 11333
rect 14836 11261 14842 11295
rect 14876 11261 14882 11295
rect 14836 11223 14882 11261
rect 14836 11189 14842 11223
rect 14876 11189 14882 11223
rect 14836 11151 14882 11189
rect 14836 11117 14842 11151
rect 14876 11117 14882 11151
rect 14836 11092 14882 11117
rect 14924 12951 14970 12954
rect 14924 12917 14930 12951
rect 14964 12917 14970 12951
rect 14924 12879 14970 12917
rect 14924 12845 14930 12879
rect 14964 12845 14970 12879
rect 14924 12807 14970 12845
rect 14924 12773 14930 12807
rect 14964 12773 14970 12807
rect 14924 12735 14970 12773
rect 14924 12701 14930 12735
rect 14964 12701 14970 12735
rect 14924 12663 14970 12701
rect 14924 12629 14930 12663
rect 14964 12629 14970 12663
rect 14924 12591 14970 12629
rect 14924 12557 14930 12591
rect 14964 12557 14970 12591
rect 14924 12519 14970 12557
rect 14924 12485 14930 12519
rect 14964 12485 14970 12519
rect 14924 12447 14970 12485
rect 14924 12413 14930 12447
rect 14964 12413 14970 12447
rect 14924 12375 14970 12413
rect 14924 12341 14930 12375
rect 14964 12341 14970 12375
rect 14924 12303 14970 12341
rect 14924 12269 14930 12303
rect 14964 12269 14970 12303
rect 14924 12231 14970 12269
rect 14924 12197 14930 12231
rect 14964 12197 14970 12231
rect 14924 12159 14970 12197
rect 14924 12125 14930 12159
rect 14964 12125 14970 12159
rect 14924 12087 14970 12125
rect 14924 12053 14930 12087
rect 14964 12053 14970 12087
rect 14924 12015 14970 12053
rect 14924 11981 14930 12015
rect 14964 11981 14970 12015
rect 14924 11943 14970 11981
rect 14924 11909 14930 11943
rect 14964 11909 14970 11943
rect 14924 11871 14970 11909
rect 14924 11837 14930 11871
rect 14964 11837 14970 11871
rect 14924 11799 14970 11837
rect 14924 11765 14930 11799
rect 14964 11765 14970 11799
rect 14924 11727 14970 11765
rect 14924 11693 14930 11727
rect 14964 11693 14970 11727
rect 14924 11655 14970 11693
rect 14924 11621 14930 11655
rect 14964 11621 14970 11655
rect 14924 11583 14970 11621
rect 14924 11549 14930 11583
rect 14964 11549 14970 11583
rect 14924 11511 14970 11549
rect 14924 11477 14930 11511
rect 14964 11477 14970 11511
rect 14924 11439 14970 11477
rect 14924 11405 14930 11439
rect 14964 11405 14970 11439
rect 14924 11367 14970 11405
rect 14924 11333 14930 11367
rect 14964 11333 14970 11367
rect 14924 11295 14970 11333
rect 14924 11261 14930 11295
rect 14964 11261 14970 11295
rect 14924 11223 14970 11261
rect 14924 11189 14930 11223
rect 14964 11189 14970 11223
rect 14924 11151 14970 11189
rect 14924 11117 14930 11151
rect 14964 11117 14970 11151
rect 14836 11070 14883 11092
rect 14924 11070 14970 11117
rect 15012 12951 15058 12989
rect 15091 13038 15156 13070
rect 15091 12986 15098 13038
rect 15150 12986 15156 13038
rect 15091 12956 15156 12986
rect 15188 13044 15237 13070
rect 15276 13068 15322 13070
rect 15188 13023 15234 13044
rect 15188 12989 15194 13023
rect 15228 12989 15234 13023
rect 15012 12917 15018 12951
rect 15052 12917 15058 12951
rect 15012 12879 15058 12917
rect 15012 12845 15018 12879
rect 15052 12845 15058 12879
rect 15012 12807 15058 12845
rect 15012 12773 15018 12807
rect 15052 12773 15058 12807
rect 15012 12735 15058 12773
rect 15012 12701 15018 12735
rect 15052 12701 15058 12735
rect 15012 12663 15058 12701
rect 15012 12629 15018 12663
rect 15052 12629 15058 12663
rect 15012 12591 15058 12629
rect 15012 12557 15018 12591
rect 15052 12557 15058 12591
rect 15012 12519 15058 12557
rect 15012 12485 15018 12519
rect 15052 12485 15058 12519
rect 15012 12447 15058 12485
rect 15012 12413 15018 12447
rect 15052 12413 15058 12447
rect 15012 12375 15058 12413
rect 15012 12341 15018 12375
rect 15052 12341 15058 12375
rect 15012 12303 15058 12341
rect 15012 12269 15018 12303
rect 15052 12269 15058 12303
rect 15012 12231 15058 12269
rect 15012 12197 15018 12231
rect 15052 12197 15058 12231
rect 15012 12159 15058 12197
rect 15012 12125 15018 12159
rect 15052 12125 15058 12159
rect 15012 12087 15058 12125
rect 15012 12053 15018 12087
rect 15052 12053 15058 12087
rect 15012 12015 15058 12053
rect 15012 11981 15018 12015
rect 15052 11981 15058 12015
rect 15012 11943 15058 11981
rect 15012 11909 15018 11943
rect 15052 11909 15058 11943
rect 15012 11871 15058 11909
rect 15012 11837 15018 11871
rect 15052 11837 15058 11871
rect 15012 11799 15058 11837
rect 15012 11765 15018 11799
rect 15052 11765 15058 11799
rect 15012 11727 15058 11765
rect 15012 11693 15018 11727
rect 15052 11693 15058 11727
rect 15012 11655 15058 11693
rect 15012 11621 15018 11655
rect 15052 11621 15058 11655
rect 15012 11583 15058 11621
rect 15012 11549 15018 11583
rect 15052 11549 15058 11583
rect 15012 11511 15058 11549
rect 15012 11477 15018 11511
rect 15052 11477 15058 11511
rect 15012 11439 15058 11477
rect 15012 11405 15018 11439
rect 15052 11405 15058 11439
rect 15012 11367 15058 11405
rect 15012 11333 15018 11367
rect 15052 11333 15058 11367
rect 15012 11295 15058 11333
rect 15012 11261 15018 11295
rect 15052 11261 15058 11295
rect 15012 11223 15058 11261
rect 15012 11189 15018 11223
rect 15052 11189 15058 11223
rect 15012 11151 15058 11189
rect 15012 11117 15018 11151
rect 15052 11117 15058 11151
rect 14659 10994 14705 11070
rect 14132 10924 14353 10970
rect 14482 10924 14705 10994
rect 14837 10970 14883 11070
rect 15012 10970 15058 11117
rect 15100 12951 15146 12956
rect 15100 12917 15106 12951
rect 15140 12917 15146 12951
rect 15100 12879 15146 12917
rect 15100 12845 15106 12879
rect 15140 12845 15146 12879
rect 15100 12807 15146 12845
rect 15100 12773 15106 12807
rect 15140 12773 15146 12807
rect 15100 12735 15146 12773
rect 15100 12701 15106 12735
rect 15140 12701 15146 12735
rect 15100 12663 15146 12701
rect 15100 12629 15106 12663
rect 15140 12629 15146 12663
rect 15100 12591 15146 12629
rect 15100 12557 15106 12591
rect 15140 12557 15146 12591
rect 15100 12519 15146 12557
rect 15100 12485 15106 12519
rect 15140 12485 15146 12519
rect 15100 12447 15146 12485
rect 15100 12413 15106 12447
rect 15140 12413 15146 12447
rect 15100 12375 15146 12413
rect 15100 12341 15106 12375
rect 15140 12341 15146 12375
rect 15100 12303 15146 12341
rect 15100 12269 15106 12303
rect 15140 12269 15146 12303
rect 15100 12231 15146 12269
rect 15100 12197 15106 12231
rect 15140 12197 15146 12231
rect 15100 12159 15146 12197
rect 15100 12125 15106 12159
rect 15140 12125 15146 12159
rect 15100 12087 15146 12125
rect 15100 12053 15106 12087
rect 15140 12053 15146 12087
rect 15100 12015 15146 12053
rect 15100 11981 15106 12015
rect 15140 11981 15146 12015
rect 15100 11943 15146 11981
rect 15100 11909 15106 11943
rect 15140 11909 15146 11943
rect 15100 11871 15146 11909
rect 15100 11837 15106 11871
rect 15140 11837 15146 11871
rect 15100 11799 15146 11837
rect 15100 11765 15106 11799
rect 15140 11765 15146 11799
rect 15100 11727 15146 11765
rect 15100 11693 15106 11727
rect 15140 11693 15146 11727
rect 15100 11655 15146 11693
rect 15100 11621 15106 11655
rect 15140 11621 15146 11655
rect 15100 11583 15146 11621
rect 15100 11549 15106 11583
rect 15140 11549 15146 11583
rect 15100 11511 15146 11549
rect 15100 11477 15106 11511
rect 15140 11477 15146 11511
rect 15100 11439 15146 11477
rect 15100 11405 15106 11439
rect 15140 11405 15146 11439
rect 15100 11367 15146 11405
rect 15100 11333 15106 11367
rect 15140 11333 15146 11367
rect 15100 11295 15146 11333
rect 15100 11261 15106 11295
rect 15140 11261 15146 11295
rect 15100 11223 15146 11261
rect 15100 11189 15106 11223
rect 15140 11189 15146 11223
rect 15100 11151 15146 11189
rect 15100 11117 15106 11151
rect 15140 11117 15146 11151
rect 15100 11070 15146 11117
rect 15188 12951 15234 12989
rect 15270 13038 15332 13068
rect 15270 12986 15275 13038
rect 15327 12986 15332 13038
rect 15270 12956 15332 12986
rect 15364 13053 15412 13070
rect 15452 13065 15498 13070
rect 15364 13023 15410 13053
rect 15364 12989 15370 13023
rect 15404 12989 15410 13023
rect 15188 12917 15194 12951
rect 15228 12917 15234 12951
rect 15188 12879 15234 12917
rect 15188 12845 15194 12879
rect 15228 12845 15234 12879
rect 15188 12807 15234 12845
rect 15188 12773 15194 12807
rect 15228 12773 15234 12807
rect 15188 12735 15234 12773
rect 15188 12701 15194 12735
rect 15228 12701 15234 12735
rect 15188 12663 15234 12701
rect 15188 12629 15194 12663
rect 15228 12629 15234 12663
rect 15188 12591 15234 12629
rect 15188 12557 15194 12591
rect 15228 12557 15234 12591
rect 15188 12519 15234 12557
rect 15188 12485 15194 12519
rect 15228 12485 15234 12519
rect 15188 12447 15234 12485
rect 15188 12413 15194 12447
rect 15228 12413 15234 12447
rect 15188 12375 15234 12413
rect 15188 12341 15194 12375
rect 15228 12341 15234 12375
rect 15188 12303 15234 12341
rect 15188 12269 15194 12303
rect 15228 12269 15234 12303
rect 15188 12231 15234 12269
rect 15188 12197 15194 12231
rect 15228 12197 15234 12231
rect 15188 12159 15234 12197
rect 15188 12125 15194 12159
rect 15228 12125 15234 12159
rect 15188 12087 15234 12125
rect 15188 12053 15194 12087
rect 15228 12053 15234 12087
rect 15188 12015 15234 12053
rect 15188 11981 15194 12015
rect 15228 11981 15234 12015
rect 15188 11943 15234 11981
rect 15188 11909 15194 11943
rect 15228 11909 15234 11943
rect 15188 11871 15234 11909
rect 15188 11837 15194 11871
rect 15228 11837 15234 11871
rect 15188 11799 15234 11837
rect 15188 11765 15194 11799
rect 15228 11765 15234 11799
rect 15188 11727 15234 11765
rect 15188 11693 15194 11727
rect 15228 11693 15234 11727
rect 15188 11655 15234 11693
rect 15188 11621 15194 11655
rect 15228 11621 15234 11655
rect 15188 11583 15234 11621
rect 15188 11549 15194 11583
rect 15228 11549 15234 11583
rect 15188 11511 15234 11549
rect 15188 11477 15194 11511
rect 15228 11477 15234 11511
rect 15188 11439 15234 11477
rect 15188 11405 15194 11439
rect 15228 11405 15234 11439
rect 15188 11367 15234 11405
rect 15188 11333 15194 11367
rect 15228 11333 15234 11367
rect 15188 11295 15234 11333
rect 15188 11261 15194 11295
rect 15228 11261 15234 11295
rect 15188 11223 15234 11261
rect 15188 11189 15194 11223
rect 15228 11189 15234 11223
rect 15188 11151 15234 11189
rect 15188 11117 15194 11151
rect 15228 11117 15234 11151
rect 15188 11092 15234 11117
rect 15276 12951 15322 12956
rect 15276 12917 15282 12951
rect 15316 12917 15322 12951
rect 15276 12879 15322 12917
rect 15276 12845 15282 12879
rect 15316 12845 15322 12879
rect 15276 12807 15322 12845
rect 15276 12773 15282 12807
rect 15316 12773 15322 12807
rect 15276 12735 15322 12773
rect 15276 12701 15282 12735
rect 15316 12701 15322 12735
rect 15276 12663 15322 12701
rect 15276 12629 15282 12663
rect 15316 12629 15322 12663
rect 15276 12591 15322 12629
rect 15276 12557 15282 12591
rect 15316 12557 15322 12591
rect 15276 12519 15322 12557
rect 15276 12485 15282 12519
rect 15316 12485 15322 12519
rect 15276 12447 15322 12485
rect 15276 12413 15282 12447
rect 15316 12413 15322 12447
rect 15276 12375 15322 12413
rect 15276 12341 15282 12375
rect 15316 12341 15322 12375
rect 15276 12303 15322 12341
rect 15276 12269 15282 12303
rect 15316 12269 15322 12303
rect 15276 12231 15322 12269
rect 15276 12197 15282 12231
rect 15316 12197 15322 12231
rect 15276 12159 15322 12197
rect 15276 12125 15282 12159
rect 15316 12125 15322 12159
rect 15276 12087 15322 12125
rect 15276 12053 15282 12087
rect 15316 12053 15322 12087
rect 15276 12015 15322 12053
rect 15276 11981 15282 12015
rect 15316 11981 15322 12015
rect 15276 11943 15322 11981
rect 15276 11909 15282 11943
rect 15316 11909 15322 11943
rect 15276 11871 15322 11909
rect 15276 11837 15282 11871
rect 15316 11837 15322 11871
rect 15276 11799 15322 11837
rect 15276 11765 15282 11799
rect 15316 11765 15322 11799
rect 15276 11727 15322 11765
rect 15276 11693 15282 11727
rect 15316 11693 15322 11727
rect 15276 11655 15322 11693
rect 15276 11621 15282 11655
rect 15316 11621 15322 11655
rect 15276 11583 15322 11621
rect 15276 11549 15282 11583
rect 15316 11549 15322 11583
rect 15276 11511 15322 11549
rect 15276 11477 15282 11511
rect 15316 11477 15322 11511
rect 15276 11439 15322 11477
rect 15276 11405 15282 11439
rect 15316 11405 15322 11439
rect 15276 11367 15322 11405
rect 15276 11333 15282 11367
rect 15316 11333 15322 11367
rect 15276 11295 15322 11333
rect 15276 11261 15282 11295
rect 15316 11261 15322 11295
rect 15276 11223 15322 11261
rect 15276 11189 15282 11223
rect 15316 11189 15322 11223
rect 15276 11151 15322 11189
rect 15276 11117 15282 11151
rect 15316 11117 15322 11151
rect 15188 11070 15236 11092
rect 15276 11070 15322 11117
rect 15364 12951 15410 12989
rect 15443 13033 15508 13065
rect 15443 12981 15450 13033
rect 15502 12981 15508 13033
rect 15443 12951 15508 12981
rect 15540 13044 15587 13070
rect 15628 13068 15674 13070
rect 15540 13023 15586 13044
rect 15540 12989 15546 13023
rect 15580 12989 15586 13023
rect 15540 12951 15586 12989
rect 15622 13038 15684 13068
rect 15622 12986 15627 13038
rect 15679 12986 15684 13038
rect 15622 12956 15684 12986
rect 15716 13051 15766 13070
rect 15804 13065 15850 13070
rect 15716 13023 15762 13051
rect 15716 12989 15722 13023
rect 15756 12989 15762 13023
rect 15364 12917 15370 12951
rect 15404 12917 15410 12951
rect 15364 12879 15410 12917
rect 15364 12845 15370 12879
rect 15404 12845 15410 12879
rect 15364 12807 15410 12845
rect 15364 12773 15370 12807
rect 15404 12773 15410 12807
rect 15364 12735 15410 12773
rect 15364 12701 15370 12735
rect 15404 12701 15410 12735
rect 15364 12663 15410 12701
rect 15364 12629 15370 12663
rect 15404 12629 15410 12663
rect 15364 12591 15410 12629
rect 15364 12557 15370 12591
rect 15404 12557 15410 12591
rect 15364 12519 15410 12557
rect 15364 12485 15370 12519
rect 15404 12485 15410 12519
rect 15364 12447 15410 12485
rect 15364 12413 15370 12447
rect 15404 12413 15410 12447
rect 15364 12375 15410 12413
rect 15364 12341 15370 12375
rect 15404 12341 15410 12375
rect 15364 12303 15410 12341
rect 15364 12269 15370 12303
rect 15404 12269 15410 12303
rect 15364 12231 15410 12269
rect 15364 12197 15370 12231
rect 15404 12197 15410 12231
rect 15364 12159 15410 12197
rect 15364 12125 15370 12159
rect 15404 12125 15410 12159
rect 15364 12087 15410 12125
rect 15364 12053 15370 12087
rect 15404 12053 15410 12087
rect 15364 12015 15410 12053
rect 15364 11981 15370 12015
rect 15404 11981 15410 12015
rect 15364 11943 15410 11981
rect 15364 11909 15370 11943
rect 15404 11909 15410 11943
rect 15364 11871 15410 11909
rect 15364 11837 15370 11871
rect 15404 11837 15410 11871
rect 15364 11799 15410 11837
rect 15364 11765 15370 11799
rect 15404 11765 15410 11799
rect 15364 11727 15410 11765
rect 15364 11693 15370 11727
rect 15404 11693 15410 11727
rect 15364 11655 15410 11693
rect 15364 11621 15370 11655
rect 15404 11621 15410 11655
rect 15364 11583 15410 11621
rect 15364 11549 15370 11583
rect 15404 11549 15410 11583
rect 15364 11511 15410 11549
rect 15364 11477 15370 11511
rect 15404 11477 15410 11511
rect 15364 11439 15410 11477
rect 15364 11405 15370 11439
rect 15404 11405 15410 11439
rect 15364 11367 15410 11405
rect 15364 11333 15370 11367
rect 15404 11333 15410 11367
rect 15364 11295 15410 11333
rect 15364 11261 15370 11295
rect 15404 11261 15410 11295
rect 15364 11223 15410 11261
rect 15364 11189 15370 11223
rect 15404 11189 15410 11223
rect 15364 11151 15410 11189
rect 15364 11117 15370 11151
rect 15404 11117 15410 11151
rect 15364 11101 15410 11117
rect 15452 12917 15458 12951
rect 15492 12917 15498 12951
rect 15452 12879 15498 12917
rect 15452 12845 15458 12879
rect 15492 12845 15498 12879
rect 15452 12807 15498 12845
rect 15452 12773 15458 12807
rect 15492 12773 15498 12807
rect 15452 12735 15498 12773
rect 15452 12701 15458 12735
rect 15492 12701 15498 12735
rect 15452 12663 15498 12701
rect 15452 12629 15458 12663
rect 15492 12629 15498 12663
rect 15452 12591 15498 12629
rect 15452 12557 15458 12591
rect 15492 12557 15498 12591
rect 15452 12519 15498 12557
rect 15452 12485 15458 12519
rect 15492 12485 15498 12519
rect 15452 12447 15498 12485
rect 15452 12413 15458 12447
rect 15492 12413 15498 12447
rect 15452 12375 15498 12413
rect 15452 12341 15458 12375
rect 15492 12341 15498 12375
rect 15452 12303 15498 12341
rect 15452 12269 15458 12303
rect 15492 12269 15498 12303
rect 15452 12231 15498 12269
rect 15452 12197 15458 12231
rect 15492 12197 15498 12231
rect 15452 12159 15498 12197
rect 15452 12125 15458 12159
rect 15492 12125 15498 12159
rect 15452 12087 15498 12125
rect 15452 12053 15458 12087
rect 15492 12053 15498 12087
rect 15452 12015 15498 12053
rect 15452 11981 15458 12015
rect 15492 11981 15498 12015
rect 15452 11943 15498 11981
rect 15452 11909 15458 11943
rect 15492 11909 15498 11943
rect 15452 11871 15498 11909
rect 15452 11837 15458 11871
rect 15492 11837 15498 11871
rect 15452 11799 15498 11837
rect 15452 11765 15458 11799
rect 15492 11765 15498 11799
rect 15452 11727 15498 11765
rect 15452 11693 15458 11727
rect 15492 11693 15498 11727
rect 15452 11655 15498 11693
rect 15452 11621 15458 11655
rect 15492 11621 15498 11655
rect 15452 11583 15498 11621
rect 15452 11549 15458 11583
rect 15492 11549 15498 11583
rect 15452 11511 15498 11549
rect 15452 11477 15458 11511
rect 15492 11477 15498 11511
rect 15452 11439 15498 11477
rect 15452 11405 15458 11439
rect 15492 11405 15498 11439
rect 15452 11367 15498 11405
rect 15452 11333 15458 11367
rect 15492 11333 15498 11367
rect 15452 11295 15498 11333
rect 15452 11261 15458 11295
rect 15492 11261 15498 11295
rect 15452 11223 15498 11261
rect 15452 11189 15458 11223
rect 15492 11189 15498 11223
rect 15452 11151 15498 11189
rect 15452 11117 15458 11151
rect 15492 11117 15498 11151
rect 15364 11070 15411 11101
rect 15452 11070 15498 11117
rect 15540 12917 15546 12951
rect 15580 12917 15586 12951
rect 15540 12879 15586 12917
rect 15540 12845 15546 12879
rect 15580 12845 15586 12879
rect 15540 12807 15586 12845
rect 15540 12773 15546 12807
rect 15580 12773 15586 12807
rect 15540 12735 15586 12773
rect 15540 12701 15546 12735
rect 15580 12701 15586 12735
rect 15540 12663 15586 12701
rect 15540 12629 15546 12663
rect 15580 12629 15586 12663
rect 15540 12591 15586 12629
rect 15540 12557 15546 12591
rect 15580 12557 15586 12591
rect 15540 12519 15586 12557
rect 15540 12485 15546 12519
rect 15580 12485 15586 12519
rect 15540 12447 15586 12485
rect 15540 12413 15546 12447
rect 15580 12413 15586 12447
rect 15540 12375 15586 12413
rect 15540 12341 15546 12375
rect 15580 12341 15586 12375
rect 15540 12303 15586 12341
rect 15540 12269 15546 12303
rect 15580 12269 15586 12303
rect 15540 12231 15586 12269
rect 15540 12197 15546 12231
rect 15580 12197 15586 12231
rect 15540 12159 15586 12197
rect 15540 12125 15546 12159
rect 15580 12125 15586 12159
rect 15540 12087 15586 12125
rect 15540 12053 15546 12087
rect 15580 12053 15586 12087
rect 15540 12015 15586 12053
rect 15540 11981 15546 12015
rect 15580 11981 15586 12015
rect 15540 11943 15586 11981
rect 15540 11909 15546 11943
rect 15580 11909 15586 11943
rect 15540 11871 15586 11909
rect 15540 11837 15546 11871
rect 15580 11837 15586 11871
rect 15540 11799 15586 11837
rect 15540 11765 15546 11799
rect 15580 11765 15586 11799
rect 15540 11727 15586 11765
rect 15540 11693 15546 11727
rect 15580 11693 15586 11727
rect 15540 11655 15586 11693
rect 15540 11621 15546 11655
rect 15580 11621 15586 11655
rect 15540 11583 15586 11621
rect 15540 11549 15546 11583
rect 15580 11549 15586 11583
rect 15540 11511 15586 11549
rect 15540 11477 15546 11511
rect 15580 11477 15586 11511
rect 15540 11439 15586 11477
rect 15540 11405 15546 11439
rect 15580 11405 15586 11439
rect 15540 11367 15586 11405
rect 15540 11333 15546 11367
rect 15580 11333 15586 11367
rect 15540 11295 15586 11333
rect 15540 11261 15546 11295
rect 15580 11261 15586 11295
rect 15540 11223 15586 11261
rect 15540 11189 15546 11223
rect 15580 11189 15586 11223
rect 15540 11151 15586 11189
rect 15540 11117 15546 11151
rect 15580 11117 15586 11151
rect 14837 10924 15058 10970
rect 15190 10970 15236 11070
rect 15365 10970 15411 11070
rect 15190 10924 15411 10970
rect 15540 10971 15586 11117
rect 15628 12951 15674 12956
rect 15628 12917 15634 12951
rect 15668 12917 15674 12951
rect 15628 12879 15674 12917
rect 15628 12845 15634 12879
rect 15668 12845 15674 12879
rect 15628 12807 15674 12845
rect 15628 12773 15634 12807
rect 15668 12773 15674 12807
rect 15628 12735 15674 12773
rect 15628 12701 15634 12735
rect 15668 12701 15674 12735
rect 15628 12663 15674 12701
rect 15628 12629 15634 12663
rect 15668 12629 15674 12663
rect 15628 12591 15674 12629
rect 15628 12557 15634 12591
rect 15668 12557 15674 12591
rect 15628 12519 15674 12557
rect 15628 12485 15634 12519
rect 15668 12485 15674 12519
rect 15628 12447 15674 12485
rect 15628 12413 15634 12447
rect 15668 12413 15674 12447
rect 15628 12375 15674 12413
rect 15628 12341 15634 12375
rect 15668 12341 15674 12375
rect 15628 12303 15674 12341
rect 15628 12269 15634 12303
rect 15668 12269 15674 12303
rect 15628 12231 15674 12269
rect 15628 12197 15634 12231
rect 15668 12197 15674 12231
rect 15628 12159 15674 12197
rect 15628 12125 15634 12159
rect 15668 12125 15674 12159
rect 15628 12087 15674 12125
rect 15628 12053 15634 12087
rect 15668 12053 15674 12087
rect 15628 12015 15674 12053
rect 15628 11981 15634 12015
rect 15668 11981 15674 12015
rect 15628 11943 15674 11981
rect 15628 11909 15634 11943
rect 15668 11909 15674 11943
rect 15628 11871 15674 11909
rect 15628 11837 15634 11871
rect 15668 11837 15674 11871
rect 15628 11799 15674 11837
rect 15628 11765 15634 11799
rect 15668 11765 15674 11799
rect 15628 11727 15674 11765
rect 15628 11693 15634 11727
rect 15668 11693 15674 11727
rect 15628 11655 15674 11693
rect 15628 11621 15634 11655
rect 15668 11621 15674 11655
rect 15628 11583 15674 11621
rect 15628 11549 15634 11583
rect 15668 11549 15674 11583
rect 15628 11511 15674 11549
rect 15628 11477 15634 11511
rect 15668 11477 15674 11511
rect 15628 11439 15674 11477
rect 15628 11405 15634 11439
rect 15668 11405 15674 11439
rect 15628 11367 15674 11405
rect 15628 11333 15634 11367
rect 15668 11333 15674 11367
rect 15628 11295 15674 11333
rect 15628 11261 15634 11295
rect 15668 11261 15674 11295
rect 15628 11223 15674 11261
rect 15628 11189 15634 11223
rect 15668 11189 15674 11223
rect 15628 11151 15674 11189
rect 15628 11117 15634 11151
rect 15668 11117 15674 11151
rect 15628 11070 15674 11117
rect 15716 12951 15762 12989
rect 15796 13033 15861 13065
rect 15796 12981 15803 13033
rect 15855 12981 15861 13033
rect 15796 12951 15861 12981
rect 15892 13042 15941 13070
rect 15980 13064 16026 13070
rect 15892 13023 15938 13042
rect 15892 12989 15898 13023
rect 15932 12989 15938 13023
rect 15892 12951 15938 12989
rect 15972 13034 16034 13064
rect 15972 12982 15977 13034
rect 16029 12982 16034 13034
rect 15972 12952 16034 12982
rect 16068 13049 16115 13070
rect 16156 13065 16202 13070
rect 16068 13023 16114 13049
rect 16068 12989 16074 13023
rect 16108 12989 16114 13023
rect 15716 12917 15722 12951
rect 15756 12917 15762 12951
rect 15716 12879 15762 12917
rect 15716 12845 15722 12879
rect 15756 12845 15762 12879
rect 15716 12807 15762 12845
rect 15716 12773 15722 12807
rect 15756 12773 15762 12807
rect 15716 12735 15762 12773
rect 15716 12701 15722 12735
rect 15756 12701 15762 12735
rect 15716 12663 15762 12701
rect 15716 12629 15722 12663
rect 15756 12629 15762 12663
rect 15716 12591 15762 12629
rect 15716 12557 15722 12591
rect 15756 12557 15762 12591
rect 15716 12519 15762 12557
rect 15716 12485 15722 12519
rect 15756 12485 15762 12519
rect 15716 12447 15762 12485
rect 15716 12413 15722 12447
rect 15756 12413 15762 12447
rect 15716 12375 15762 12413
rect 15716 12341 15722 12375
rect 15756 12341 15762 12375
rect 15716 12303 15762 12341
rect 15716 12269 15722 12303
rect 15756 12269 15762 12303
rect 15716 12231 15762 12269
rect 15716 12197 15722 12231
rect 15756 12197 15762 12231
rect 15716 12159 15762 12197
rect 15716 12125 15722 12159
rect 15756 12125 15762 12159
rect 15716 12087 15762 12125
rect 15716 12053 15722 12087
rect 15756 12053 15762 12087
rect 15716 12015 15762 12053
rect 15716 11981 15722 12015
rect 15756 11981 15762 12015
rect 15716 11943 15762 11981
rect 15716 11909 15722 11943
rect 15756 11909 15762 11943
rect 15716 11871 15762 11909
rect 15716 11837 15722 11871
rect 15756 11837 15762 11871
rect 15716 11799 15762 11837
rect 15716 11765 15722 11799
rect 15756 11765 15762 11799
rect 15716 11727 15762 11765
rect 15716 11693 15722 11727
rect 15756 11693 15762 11727
rect 15716 11655 15762 11693
rect 15716 11621 15722 11655
rect 15756 11621 15762 11655
rect 15716 11583 15762 11621
rect 15716 11549 15722 11583
rect 15756 11549 15762 11583
rect 15716 11511 15762 11549
rect 15716 11477 15722 11511
rect 15756 11477 15762 11511
rect 15716 11439 15762 11477
rect 15716 11405 15722 11439
rect 15756 11405 15762 11439
rect 15716 11367 15762 11405
rect 15716 11333 15722 11367
rect 15756 11333 15762 11367
rect 15716 11295 15762 11333
rect 15716 11261 15722 11295
rect 15756 11261 15762 11295
rect 15716 11223 15762 11261
rect 15716 11189 15722 11223
rect 15756 11189 15762 11223
rect 15716 11151 15762 11189
rect 15716 11117 15722 11151
rect 15756 11117 15762 11151
rect 15716 11102 15762 11117
rect 15715 11070 15762 11102
rect 15804 12917 15810 12951
rect 15844 12917 15850 12951
rect 15804 12879 15850 12917
rect 15804 12845 15810 12879
rect 15844 12845 15850 12879
rect 15804 12807 15850 12845
rect 15804 12773 15810 12807
rect 15844 12773 15850 12807
rect 15804 12735 15850 12773
rect 15804 12701 15810 12735
rect 15844 12701 15850 12735
rect 15804 12663 15850 12701
rect 15804 12629 15810 12663
rect 15844 12629 15850 12663
rect 15804 12591 15850 12629
rect 15804 12557 15810 12591
rect 15844 12557 15850 12591
rect 15804 12519 15850 12557
rect 15804 12485 15810 12519
rect 15844 12485 15850 12519
rect 15804 12447 15850 12485
rect 15804 12413 15810 12447
rect 15844 12413 15850 12447
rect 15804 12375 15850 12413
rect 15804 12341 15810 12375
rect 15844 12341 15850 12375
rect 15804 12303 15850 12341
rect 15804 12269 15810 12303
rect 15844 12269 15850 12303
rect 15804 12231 15850 12269
rect 15804 12197 15810 12231
rect 15844 12197 15850 12231
rect 15804 12159 15850 12197
rect 15804 12125 15810 12159
rect 15844 12125 15850 12159
rect 15804 12087 15850 12125
rect 15804 12053 15810 12087
rect 15844 12053 15850 12087
rect 15804 12015 15850 12053
rect 15804 11981 15810 12015
rect 15844 11981 15850 12015
rect 15804 11943 15850 11981
rect 15804 11909 15810 11943
rect 15844 11909 15850 11943
rect 15804 11871 15850 11909
rect 15804 11837 15810 11871
rect 15844 11837 15850 11871
rect 15804 11799 15850 11837
rect 15804 11765 15810 11799
rect 15844 11765 15850 11799
rect 15804 11727 15850 11765
rect 15804 11693 15810 11727
rect 15844 11693 15850 11727
rect 15804 11655 15850 11693
rect 15804 11621 15810 11655
rect 15844 11621 15850 11655
rect 15804 11583 15850 11621
rect 15804 11549 15810 11583
rect 15844 11549 15850 11583
rect 15804 11511 15850 11549
rect 15804 11477 15810 11511
rect 15844 11477 15850 11511
rect 15804 11439 15850 11477
rect 15804 11405 15810 11439
rect 15844 11405 15850 11439
rect 15804 11367 15850 11405
rect 15804 11333 15810 11367
rect 15844 11333 15850 11367
rect 15804 11295 15850 11333
rect 15804 11261 15810 11295
rect 15844 11261 15850 11295
rect 15804 11223 15850 11261
rect 15804 11189 15810 11223
rect 15844 11189 15850 11223
rect 15804 11151 15850 11189
rect 15804 11117 15810 11151
rect 15844 11117 15850 11151
rect 15804 11070 15850 11117
rect 15892 12917 15898 12951
rect 15932 12917 15938 12951
rect 15892 12879 15938 12917
rect 15892 12845 15898 12879
rect 15932 12845 15938 12879
rect 15892 12807 15938 12845
rect 15892 12773 15898 12807
rect 15932 12773 15938 12807
rect 15892 12735 15938 12773
rect 15892 12701 15898 12735
rect 15932 12701 15938 12735
rect 15892 12663 15938 12701
rect 15892 12629 15898 12663
rect 15932 12629 15938 12663
rect 15892 12591 15938 12629
rect 15892 12557 15898 12591
rect 15932 12557 15938 12591
rect 15892 12519 15938 12557
rect 15892 12485 15898 12519
rect 15932 12485 15938 12519
rect 15892 12447 15938 12485
rect 15892 12413 15898 12447
rect 15932 12413 15938 12447
rect 15892 12375 15938 12413
rect 15892 12341 15898 12375
rect 15932 12341 15938 12375
rect 15892 12303 15938 12341
rect 15892 12269 15898 12303
rect 15932 12269 15938 12303
rect 15892 12231 15938 12269
rect 15892 12197 15898 12231
rect 15932 12197 15938 12231
rect 15892 12159 15938 12197
rect 15892 12125 15898 12159
rect 15932 12125 15938 12159
rect 15892 12087 15938 12125
rect 15892 12053 15898 12087
rect 15932 12053 15938 12087
rect 15892 12015 15938 12053
rect 15892 11981 15898 12015
rect 15932 11981 15938 12015
rect 15892 11943 15938 11981
rect 15892 11909 15898 11943
rect 15932 11909 15938 11943
rect 15892 11871 15938 11909
rect 15892 11837 15898 11871
rect 15932 11837 15938 11871
rect 15892 11799 15938 11837
rect 15892 11765 15898 11799
rect 15932 11765 15938 11799
rect 15892 11727 15938 11765
rect 15892 11693 15898 11727
rect 15932 11693 15938 11727
rect 15892 11655 15938 11693
rect 15892 11621 15898 11655
rect 15932 11621 15938 11655
rect 15892 11583 15938 11621
rect 15892 11549 15898 11583
rect 15932 11549 15938 11583
rect 15892 11511 15938 11549
rect 15892 11477 15898 11511
rect 15932 11477 15938 11511
rect 15892 11439 15938 11477
rect 15892 11405 15898 11439
rect 15932 11405 15938 11439
rect 15892 11367 15938 11405
rect 15892 11333 15898 11367
rect 15932 11333 15938 11367
rect 15892 11295 15938 11333
rect 15892 11261 15898 11295
rect 15932 11261 15938 11295
rect 15892 11223 15938 11261
rect 15892 11189 15898 11223
rect 15932 11189 15938 11223
rect 15892 11151 15938 11189
rect 15892 11117 15898 11151
rect 15932 11117 15938 11151
rect 15892 11093 15938 11117
rect 15980 12951 16026 12952
rect 15980 12917 15986 12951
rect 16020 12917 16026 12951
rect 15980 12879 16026 12917
rect 15980 12845 15986 12879
rect 16020 12845 16026 12879
rect 15980 12807 16026 12845
rect 15980 12773 15986 12807
rect 16020 12773 16026 12807
rect 15980 12735 16026 12773
rect 15980 12701 15986 12735
rect 16020 12701 16026 12735
rect 15980 12663 16026 12701
rect 15980 12629 15986 12663
rect 16020 12629 16026 12663
rect 15980 12591 16026 12629
rect 15980 12557 15986 12591
rect 16020 12557 16026 12591
rect 15980 12519 16026 12557
rect 15980 12485 15986 12519
rect 16020 12485 16026 12519
rect 15980 12447 16026 12485
rect 15980 12413 15986 12447
rect 16020 12413 16026 12447
rect 15980 12375 16026 12413
rect 15980 12341 15986 12375
rect 16020 12341 16026 12375
rect 15980 12303 16026 12341
rect 15980 12269 15986 12303
rect 16020 12269 16026 12303
rect 15980 12231 16026 12269
rect 15980 12197 15986 12231
rect 16020 12197 16026 12231
rect 15980 12159 16026 12197
rect 15980 12125 15986 12159
rect 16020 12125 16026 12159
rect 15980 12087 16026 12125
rect 15980 12053 15986 12087
rect 16020 12053 16026 12087
rect 15980 12015 16026 12053
rect 15980 11981 15986 12015
rect 16020 11981 16026 12015
rect 15980 11943 16026 11981
rect 15980 11909 15986 11943
rect 16020 11909 16026 11943
rect 15980 11871 16026 11909
rect 15980 11837 15986 11871
rect 16020 11837 16026 11871
rect 15980 11799 16026 11837
rect 15980 11765 15986 11799
rect 16020 11765 16026 11799
rect 15980 11727 16026 11765
rect 15980 11693 15986 11727
rect 16020 11693 16026 11727
rect 15980 11655 16026 11693
rect 15980 11621 15986 11655
rect 16020 11621 16026 11655
rect 15980 11583 16026 11621
rect 15980 11549 15986 11583
rect 16020 11549 16026 11583
rect 15980 11511 16026 11549
rect 15980 11477 15986 11511
rect 16020 11477 16026 11511
rect 15980 11439 16026 11477
rect 15980 11405 15986 11439
rect 16020 11405 16026 11439
rect 15980 11367 16026 11405
rect 15980 11333 15986 11367
rect 16020 11333 16026 11367
rect 15980 11295 16026 11333
rect 15980 11261 15986 11295
rect 16020 11261 16026 11295
rect 15980 11223 16026 11261
rect 15980 11189 15986 11223
rect 16020 11189 16026 11223
rect 15980 11151 16026 11189
rect 15980 11117 15986 11151
rect 16020 11117 16026 11151
rect 15892 11070 15941 11093
rect 15980 11070 16026 11117
rect 16068 12951 16114 12989
rect 16148 13033 16213 13065
rect 16148 12981 16155 13033
rect 16207 12981 16213 13033
rect 16148 12951 16213 12981
rect 16244 13023 16290 13171
rect 16423 13175 16644 13221
rect 16423 13070 16469 13175
rect 16598 13070 16644 13175
rect 16777 13171 16998 13217
rect 16777 13070 16823 13171
rect 16952 13070 16998 13171
rect 17130 13171 17351 13217
rect 17130 13070 17176 13171
rect 17305 13070 17351 13171
rect 16332 13064 16378 13070
rect 16244 12989 16250 13023
rect 16284 12989 16290 13023
rect 16244 12951 16290 12989
rect 16326 13034 16388 13064
rect 16326 12982 16331 13034
rect 16383 12982 16388 13034
rect 16326 12952 16388 12982
rect 16420 13053 16469 13070
rect 16508 13064 16554 13070
rect 16420 13023 16466 13053
rect 16420 12989 16426 13023
rect 16460 12989 16466 13023
rect 16068 12917 16074 12951
rect 16108 12917 16114 12951
rect 16068 12879 16114 12917
rect 16068 12845 16074 12879
rect 16108 12845 16114 12879
rect 16068 12807 16114 12845
rect 16068 12773 16074 12807
rect 16108 12773 16114 12807
rect 16068 12735 16114 12773
rect 16068 12701 16074 12735
rect 16108 12701 16114 12735
rect 16068 12663 16114 12701
rect 16068 12629 16074 12663
rect 16108 12629 16114 12663
rect 16068 12591 16114 12629
rect 16068 12557 16074 12591
rect 16108 12557 16114 12591
rect 16068 12519 16114 12557
rect 16068 12485 16074 12519
rect 16108 12485 16114 12519
rect 16068 12447 16114 12485
rect 16068 12413 16074 12447
rect 16108 12413 16114 12447
rect 16068 12375 16114 12413
rect 16068 12341 16074 12375
rect 16108 12341 16114 12375
rect 16068 12303 16114 12341
rect 16068 12269 16074 12303
rect 16108 12269 16114 12303
rect 16068 12231 16114 12269
rect 16068 12197 16074 12231
rect 16108 12197 16114 12231
rect 16068 12159 16114 12197
rect 16068 12125 16074 12159
rect 16108 12125 16114 12159
rect 16068 12087 16114 12125
rect 16068 12053 16074 12087
rect 16108 12053 16114 12087
rect 16068 12015 16114 12053
rect 16068 11981 16074 12015
rect 16108 11981 16114 12015
rect 16068 11943 16114 11981
rect 16068 11909 16074 11943
rect 16108 11909 16114 11943
rect 16068 11871 16114 11909
rect 16068 11837 16074 11871
rect 16108 11837 16114 11871
rect 16068 11799 16114 11837
rect 16068 11765 16074 11799
rect 16108 11765 16114 11799
rect 16068 11727 16114 11765
rect 16068 11693 16074 11727
rect 16108 11693 16114 11727
rect 16068 11655 16114 11693
rect 16068 11621 16074 11655
rect 16108 11621 16114 11655
rect 16068 11583 16114 11621
rect 16068 11549 16074 11583
rect 16108 11549 16114 11583
rect 16068 11511 16114 11549
rect 16068 11477 16074 11511
rect 16108 11477 16114 11511
rect 16068 11439 16114 11477
rect 16068 11405 16074 11439
rect 16108 11405 16114 11439
rect 16068 11367 16114 11405
rect 16068 11333 16074 11367
rect 16108 11333 16114 11367
rect 16068 11295 16114 11333
rect 16068 11261 16074 11295
rect 16108 11261 16114 11295
rect 16068 11223 16114 11261
rect 16068 11189 16074 11223
rect 16108 11189 16114 11223
rect 16068 11151 16114 11189
rect 16068 11117 16074 11151
rect 16108 11117 16114 11151
rect 16068 11102 16114 11117
rect 16156 12917 16162 12951
rect 16196 12917 16202 12951
rect 16156 12879 16202 12917
rect 16156 12845 16162 12879
rect 16196 12845 16202 12879
rect 16156 12807 16202 12845
rect 16156 12773 16162 12807
rect 16196 12773 16202 12807
rect 16156 12735 16202 12773
rect 16156 12701 16162 12735
rect 16196 12701 16202 12735
rect 16156 12663 16202 12701
rect 16156 12629 16162 12663
rect 16196 12629 16202 12663
rect 16156 12591 16202 12629
rect 16156 12557 16162 12591
rect 16196 12557 16202 12591
rect 16156 12519 16202 12557
rect 16156 12485 16162 12519
rect 16196 12485 16202 12519
rect 16156 12447 16202 12485
rect 16156 12413 16162 12447
rect 16196 12413 16202 12447
rect 16156 12375 16202 12413
rect 16156 12341 16162 12375
rect 16196 12341 16202 12375
rect 16156 12303 16202 12341
rect 16156 12269 16162 12303
rect 16196 12269 16202 12303
rect 16156 12231 16202 12269
rect 16156 12197 16162 12231
rect 16196 12197 16202 12231
rect 16156 12159 16202 12197
rect 16156 12125 16162 12159
rect 16196 12125 16202 12159
rect 16156 12087 16202 12125
rect 16156 12053 16162 12087
rect 16196 12053 16202 12087
rect 16156 12015 16202 12053
rect 16156 11981 16162 12015
rect 16196 11981 16202 12015
rect 16156 11943 16202 11981
rect 16156 11909 16162 11943
rect 16196 11909 16202 11943
rect 16156 11871 16202 11909
rect 16156 11837 16162 11871
rect 16196 11837 16202 11871
rect 16156 11799 16202 11837
rect 16156 11765 16162 11799
rect 16196 11765 16202 11799
rect 16156 11727 16202 11765
rect 16156 11693 16162 11727
rect 16196 11693 16202 11727
rect 16156 11655 16202 11693
rect 16156 11621 16162 11655
rect 16196 11621 16202 11655
rect 16156 11583 16202 11621
rect 16156 11549 16162 11583
rect 16196 11549 16202 11583
rect 16156 11511 16202 11549
rect 16156 11477 16162 11511
rect 16196 11477 16202 11511
rect 16156 11439 16202 11477
rect 16156 11405 16162 11439
rect 16196 11405 16202 11439
rect 16156 11367 16202 11405
rect 16156 11333 16162 11367
rect 16196 11333 16202 11367
rect 16156 11295 16202 11333
rect 16156 11261 16162 11295
rect 16196 11261 16202 11295
rect 16156 11223 16202 11261
rect 16156 11189 16162 11223
rect 16196 11189 16202 11223
rect 16156 11151 16202 11189
rect 16156 11117 16162 11151
rect 16196 11117 16202 11151
rect 16068 11070 16116 11102
rect 16156 11070 16202 11117
rect 16244 12917 16250 12951
rect 16284 12917 16290 12951
rect 16244 12879 16290 12917
rect 16244 12845 16250 12879
rect 16284 12845 16290 12879
rect 16244 12807 16290 12845
rect 16244 12773 16250 12807
rect 16284 12773 16290 12807
rect 16244 12735 16290 12773
rect 16244 12701 16250 12735
rect 16284 12701 16290 12735
rect 16244 12663 16290 12701
rect 16244 12629 16250 12663
rect 16284 12629 16290 12663
rect 16244 12591 16290 12629
rect 16244 12557 16250 12591
rect 16284 12557 16290 12591
rect 16244 12519 16290 12557
rect 16244 12485 16250 12519
rect 16284 12485 16290 12519
rect 16244 12447 16290 12485
rect 16244 12413 16250 12447
rect 16284 12413 16290 12447
rect 16244 12375 16290 12413
rect 16244 12341 16250 12375
rect 16284 12341 16290 12375
rect 16244 12303 16290 12341
rect 16244 12269 16250 12303
rect 16284 12269 16290 12303
rect 16244 12231 16290 12269
rect 16244 12197 16250 12231
rect 16284 12197 16290 12231
rect 16244 12159 16290 12197
rect 16244 12125 16250 12159
rect 16284 12125 16290 12159
rect 16244 12087 16290 12125
rect 16244 12053 16250 12087
rect 16284 12053 16290 12087
rect 16244 12015 16290 12053
rect 16244 11981 16250 12015
rect 16284 11981 16290 12015
rect 16244 11943 16290 11981
rect 16244 11909 16250 11943
rect 16284 11909 16290 11943
rect 16244 11871 16290 11909
rect 16244 11837 16250 11871
rect 16284 11837 16290 11871
rect 16244 11799 16290 11837
rect 16244 11765 16250 11799
rect 16284 11765 16290 11799
rect 16244 11727 16290 11765
rect 16244 11693 16250 11727
rect 16284 11693 16290 11727
rect 16244 11655 16290 11693
rect 16244 11621 16250 11655
rect 16284 11621 16290 11655
rect 16244 11583 16290 11621
rect 16244 11549 16250 11583
rect 16284 11549 16290 11583
rect 16244 11511 16290 11549
rect 16244 11477 16250 11511
rect 16284 11477 16290 11511
rect 16244 11439 16290 11477
rect 16244 11405 16250 11439
rect 16284 11405 16290 11439
rect 16244 11367 16290 11405
rect 16244 11333 16250 11367
rect 16284 11333 16290 11367
rect 16244 11295 16290 11333
rect 16244 11261 16250 11295
rect 16284 11261 16290 11295
rect 16244 11223 16290 11261
rect 16244 11189 16250 11223
rect 16284 11189 16290 11223
rect 16244 11151 16290 11189
rect 16244 11117 16250 11151
rect 16284 11117 16290 11151
rect 15715 10971 15761 11070
rect 15540 10925 15761 10971
rect 15895 10971 15941 11070
rect 16070 10971 16116 11070
rect 15895 10925 16116 10971
rect 16244 10971 16290 11117
rect 16332 12951 16378 12952
rect 16332 12917 16338 12951
rect 16372 12917 16378 12951
rect 16332 12879 16378 12917
rect 16332 12845 16338 12879
rect 16372 12845 16378 12879
rect 16332 12807 16378 12845
rect 16332 12773 16338 12807
rect 16372 12773 16378 12807
rect 16332 12735 16378 12773
rect 16332 12701 16338 12735
rect 16372 12701 16378 12735
rect 16332 12663 16378 12701
rect 16332 12629 16338 12663
rect 16372 12629 16378 12663
rect 16332 12591 16378 12629
rect 16332 12557 16338 12591
rect 16372 12557 16378 12591
rect 16332 12519 16378 12557
rect 16332 12485 16338 12519
rect 16372 12485 16378 12519
rect 16332 12447 16378 12485
rect 16332 12413 16338 12447
rect 16372 12413 16378 12447
rect 16332 12375 16378 12413
rect 16332 12341 16338 12375
rect 16372 12341 16378 12375
rect 16332 12303 16378 12341
rect 16332 12269 16338 12303
rect 16372 12269 16378 12303
rect 16332 12231 16378 12269
rect 16332 12197 16338 12231
rect 16372 12197 16378 12231
rect 16332 12159 16378 12197
rect 16332 12125 16338 12159
rect 16372 12125 16378 12159
rect 16332 12087 16378 12125
rect 16332 12053 16338 12087
rect 16372 12053 16378 12087
rect 16332 12015 16378 12053
rect 16332 11981 16338 12015
rect 16372 11981 16378 12015
rect 16332 11943 16378 11981
rect 16332 11909 16338 11943
rect 16372 11909 16378 11943
rect 16332 11871 16378 11909
rect 16332 11837 16338 11871
rect 16372 11837 16378 11871
rect 16332 11799 16378 11837
rect 16332 11765 16338 11799
rect 16372 11765 16378 11799
rect 16332 11727 16378 11765
rect 16332 11693 16338 11727
rect 16372 11693 16378 11727
rect 16332 11655 16378 11693
rect 16332 11621 16338 11655
rect 16372 11621 16378 11655
rect 16332 11583 16378 11621
rect 16332 11549 16338 11583
rect 16372 11549 16378 11583
rect 16332 11511 16378 11549
rect 16332 11477 16338 11511
rect 16372 11477 16378 11511
rect 16332 11439 16378 11477
rect 16332 11405 16338 11439
rect 16372 11405 16378 11439
rect 16332 11367 16378 11405
rect 16332 11333 16338 11367
rect 16372 11333 16378 11367
rect 16332 11295 16378 11333
rect 16332 11261 16338 11295
rect 16372 11261 16378 11295
rect 16332 11223 16378 11261
rect 16332 11189 16338 11223
rect 16372 11189 16378 11223
rect 16332 11151 16378 11189
rect 16332 11117 16338 11151
rect 16372 11117 16378 11151
rect 16332 11070 16378 11117
rect 16420 12951 16466 12989
rect 16420 12917 16426 12951
rect 16460 12917 16466 12951
rect 16502 13032 16567 13064
rect 16502 12980 16509 13032
rect 16561 12980 16567 13032
rect 16502 12951 16567 12980
rect 16502 12950 16514 12951
rect 16420 12879 16466 12917
rect 16420 12845 16426 12879
rect 16460 12845 16466 12879
rect 16420 12807 16466 12845
rect 16420 12773 16426 12807
rect 16460 12773 16466 12807
rect 16420 12735 16466 12773
rect 16420 12701 16426 12735
rect 16460 12701 16466 12735
rect 16420 12663 16466 12701
rect 16420 12629 16426 12663
rect 16460 12629 16466 12663
rect 16420 12591 16466 12629
rect 16420 12557 16426 12591
rect 16460 12557 16466 12591
rect 16420 12519 16466 12557
rect 16420 12485 16426 12519
rect 16460 12485 16466 12519
rect 16420 12447 16466 12485
rect 16420 12413 16426 12447
rect 16460 12413 16466 12447
rect 16420 12375 16466 12413
rect 16420 12341 16426 12375
rect 16460 12341 16466 12375
rect 16420 12303 16466 12341
rect 16420 12269 16426 12303
rect 16460 12269 16466 12303
rect 16420 12231 16466 12269
rect 16420 12197 16426 12231
rect 16460 12197 16466 12231
rect 16420 12159 16466 12197
rect 16420 12125 16426 12159
rect 16460 12125 16466 12159
rect 16420 12087 16466 12125
rect 16420 12053 16426 12087
rect 16460 12053 16466 12087
rect 16420 12015 16466 12053
rect 16420 11981 16426 12015
rect 16460 11981 16466 12015
rect 16420 11943 16466 11981
rect 16420 11909 16426 11943
rect 16460 11909 16466 11943
rect 16420 11871 16466 11909
rect 16420 11837 16426 11871
rect 16460 11837 16466 11871
rect 16420 11799 16466 11837
rect 16420 11765 16426 11799
rect 16460 11765 16466 11799
rect 16420 11727 16466 11765
rect 16420 11693 16426 11727
rect 16460 11693 16466 11727
rect 16420 11655 16466 11693
rect 16420 11621 16426 11655
rect 16460 11621 16466 11655
rect 16420 11583 16466 11621
rect 16420 11549 16426 11583
rect 16460 11549 16466 11583
rect 16420 11511 16466 11549
rect 16420 11477 16426 11511
rect 16460 11477 16466 11511
rect 16420 11439 16466 11477
rect 16420 11405 16426 11439
rect 16460 11405 16466 11439
rect 16420 11367 16466 11405
rect 16420 11333 16426 11367
rect 16460 11333 16466 11367
rect 16420 11295 16466 11333
rect 16420 11261 16426 11295
rect 16460 11261 16466 11295
rect 16420 11223 16466 11261
rect 16420 11189 16426 11223
rect 16460 11189 16466 11223
rect 16420 11151 16466 11189
rect 16420 11117 16426 11151
rect 16460 11117 16466 11151
rect 16420 11102 16466 11117
rect 16419 11070 16466 11102
rect 16508 12917 16514 12950
rect 16548 12950 16567 12951
rect 16596 13044 16644 13070
rect 16684 13066 16730 13070
rect 16596 13023 16642 13044
rect 16596 12989 16602 13023
rect 16636 12989 16642 13023
rect 16596 12951 16642 12989
rect 16676 13036 16738 13066
rect 16676 12984 16681 13036
rect 16733 12984 16738 13036
rect 16676 12954 16738 12984
rect 16772 13049 16823 13070
rect 16772 13023 16818 13049
rect 16772 12989 16778 13023
rect 16812 12989 16818 13023
rect 16548 12917 16554 12950
rect 16508 12879 16554 12917
rect 16508 12845 16514 12879
rect 16548 12845 16554 12879
rect 16508 12807 16554 12845
rect 16508 12773 16514 12807
rect 16548 12773 16554 12807
rect 16508 12735 16554 12773
rect 16508 12701 16514 12735
rect 16548 12701 16554 12735
rect 16508 12663 16554 12701
rect 16508 12629 16514 12663
rect 16548 12629 16554 12663
rect 16508 12591 16554 12629
rect 16508 12557 16514 12591
rect 16548 12557 16554 12591
rect 16508 12519 16554 12557
rect 16508 12485 16514 12519
rect 16548 12485 16554 12519
rect 16508 12447 16554 12485
rect 16508 12413 16514 12447
rect 16548 12413 16554 12447
rect 16508 12375 16554 12413
rect 16508 12341 16514 12375
rect 16548 12341 16554 12375
rect 16508 12303 16554 12341
rect 16508 12269 16514 12303
rect 16548 12269 16554 12303
rect 16508 12231 16554 12269
rect 16508 12197 16514 12231
rect 16548 12197 16554 12231
rect 16508 12159 16554 12197
rect 16508 12125 16514 12159
rect 16548 12125 16554 12159
rect 16508 12087 16554 12125
rect 16508 12053 16514 12087
rect 16548 12053 16554 12087
rect 16508 12015 16554 12053
rect 16508 11981 16514 12015
rect 16548 11981 16554 12015
rect 16508 11943 16554 11981
rect 16508 11909 16514 11943
rect 16548 11909 16554 11943
rect 16508 11871 16554 11909
rect 16508 11837 16514 11871
rect 16548 11837 16554 11871
rect 16508 11799 16554 11837
rect 16508 11765 16514 11799
rect 16548 11765 16554 11799
rect 16508 11727 16554 11765
rect 16508 11693 16514 11727
rect 16548 11693 16554 11727
rect 16508 11655 16554 11693
rect 16508 11621 16514 11655
rect 16548 11621 16554 11655
rect 16508 11583 16554 11621
rect 16508 11549 16514 11583
rect 16548 11549 16554 11583
rect 16508 11511 16554 11549
rect 16508 11477 16514 11511
rect 16548 11477 16554 11511
rect 16508 11439 16554 11477
rect 16508 11405 16514 11439
rect 16548 11405 16554 11439
rect 16508 11367 16554 11405
rect 16508 11333 16514 11367
rect 16548 11333 16554 11367
rect 16508 11295 16554 11333
rect 16508 11261 16514 11295
rect 16548 11261 16554 11295
rect 16508 11223 16554 11261
rect 16508 11189 16514 11223
rect 16548 11189 16554 11223
rect 16508 11151 16554 11189
rect 16508 11117 16514 11151
rect 16548 11117 16554 11151
rect 16508 11070 16554 11117
rect 16596 12917 16602 12951
rect 16636 12917 16642 12951
rect 16596 12879 16642 12917
rect 16596 12845 16602 12879
rect 16636 12845 16642 12879
rect 16596 12807 16642 12845
rect 16596 12773 16602 12807
rect 16636 12773 16642 12807
rect 16596 12735 16642 12773
rect 16596 12701 16602 12735
rect 16636 12701 16642 12735
rect 16596 12663 16642 12701
rect 16596 12629 16602 12663
rect 16636 12629 16642 12663
rect 16596 12591 16642 12629
rect 16596 12557 16602 12591
rect 16636 12557 16642 12591
rect 16596 12519 16642 12557
rect 16596 12485 16602 12519
rect 16636 12485 16642 12519
rect 16596 12447 16642 12485
rect 16596 12413 16602 12447
rect 16636 12413 16642 12447
rect 16596 12375 16642 12413
rect 16596 12341 16602 12375
rect 16636 12341 16642 12375
rect 16596 12303 16642 12341
rect 16596 12269 16602 12303
rect 16636 12269 16642 12303
rect 16596 12231 16642 12269
rect 16596 12197 16602 12231
rect 16636 12197 16642 12231
rect 16596 12159 16642 12197
rect 16596 12125 16602 12159
rect 16636 12125 16642 12159
rect 16596 12087 16642 12125
rect 16596 12053 16602 12087
rect 16636 12053 16642 12087
rect 16596 12015 16642 12053
rect 16596 11981 16602 12015
rect 16636 11981 16642 12015
rect 16596 11943 16642 11981
rect 16596 11909 16602 11943
rect 16636 11909 16642 11943
rect 16596 11871 16642 11909
rect 16596 11837 16602 11871
rect 16636 11837 16642 11871
rect 16596 11799 16642 11837
rect 16596 11765 16602 11799
rect 16636 11765 16642 11799
rect 16596 11727 16642 11765
rect 16596 11693 16602 11727
rect 16636 11693 16642 11727
rect 16596 11655 16642 11693
rect 16596 11621 16602 11655
rect 16636 11621 16642 11655
rect 16596 11583 16642 11621
rect 16596 11549 16602 11583
rect 16636 11549 16642 11583
rect 16596 11511 16642 11549
rect 16596 11477 16602 11511
rect 16636 11477 16642 11511
rect 16596 11439 16642 11477
rect 16596 11405 16602 11439
rect 16636 11405 16642 11439
rect 16596 11367 16642 11405
rect 16596 11333 16602 11367
rect 16636 11333 16642 11367
rect 16596 11295 16642 11333
rect 16596 11261 16602 11295
rect 16636 11261 16642 11295
rect 16596 11223 16642 11261
rect 16596 11189 16602 11223
rect 16636 11189 16642 11223
rect 16596 11151 16642 11189
rect 16596 11117 16602 11151
rect 16636 11117 16642 11151
rect 16419 10971 16465 11070
rect 16244 10925 16465 10971
rect 16596 10970 16642 11117
rect 16684 12951 16730 12954
rect 16684 12917 16690 12951
rect 16724 12917 16730 12951
rect 16684 12879 16730 12917
rect 16684 12845 16690 12879
rect 16724 12845 16730 12879
rect 16684 12807 16730 12845
rect 16684 12773 16690 12807
rect 16724 12773 16730 12807
rect 16684 12735 16730 12773
rect 16684 12701 16690 12735
rect 16724 12701 16730 12735
rect 16684 12663 16730 12701
rect 16684 12629 16690 12663
rect 16724 12629 16730 12663
rect 16684 12591 16730 12629
rect 16684 12557 16690 12591
rect 16724 12557 16730 12591
rect 16684 12519 16730 12557
rect 16684 12485 16690 12519
rect 16724 12485 16730 12519
rect 16684 12447 16730 12485
rect 16684 12413 16690 12447
rect 16724 12413 16730 12447
rect 16684 12375 16730 12413
rect 16684 12341 16690 12375
rect 16724 12341 16730 12375
rect 16684 12303 16730 12341
rect 16684 12269 16690 12303
rect 16724 12269 16730 12303
rect 16684 12231 16730 12269
rect 16684 12197 16690 12231
rect 16724 12197 16730 12231
rect 16684 12159 16730 12197
rect 16684 12125 16690 12159
rect 16724 12125 16730 12159
rect 16684 12087 16730 12125
rect 16684 12053 16690 12087
rect 16724 12053 16730 12087
rect 16684 12015 16730 12053
rect 16684 11981 16690 12015
rect 16724 11981 16730 12015
rect 16684 11943 16730 11981
rect 16684 11909 16690 11943
rect 16724 11909 16730 11943
rect 16684 11871 16730 11909
rect 16684 11837 16690 11871
rect 16724 11837 16730 11871
rect 16684 11799 16730 11837
rect 16684 11765 16690 11799
rect 16724 11765 16730 11799
rect 16684 11727 16730 11765
rect 16684 11693 16690 11727
rect 16724 11693 16730 11727
rect 16684 11655 16730 11693
rect 16684 11621 16690 11655
rect 16724 11621 16730 11655
rect 16684 11583 16730 11621
rect 16684 11549 16690 11583
rect 16724 11549 16730 11583
rect 16684 11511 16730 11549
rect 16684 11477 16690 11511
rect 16724 11477 16730 11511
rect 16684 11439 16730 11477
rect 16684 11405 16690 11439
rect 16724 11405 16730 11439
rect 16684 11367 16730 11405
rect 16684 11333 16690 11367
rect 16724 11333 16730 11367
rect 16684 11295 16730 11333
rect 16684 11261 16690 11295
rect 16724 11261 16730 11295
rect 16684 11223 16730 11261
rect 16684 11189 16690 11223
rect 16724 11189 16730 11223
rect 16684 11151 16730 11189
rect 16684 11117 16690 11151
rect 16724 11117 16730 11151
rect 16684 11070 16730 11117
rect 16772 12951 16818 12989
rect 16851 13038 16916 13070
rect 16851 12986 16858 13038
rect 16910 12986 16916 13038
rect 16851 12956 16916 12986
rect 16948 13040 16998 13070
rect 17036 13066 17082 13070
rect 16948 13023 16994 13040
rect 16948 12989 16954 13023
rect 16988 12989 16994 13023
rect 16772 12917 16778 12951
rect 16812 12917 16818 12951
rect 16772 12879 16818 12917
rect 16772 12845 16778 12879
rect 16812 12845 16818 12879
rect 16772 12807 16818 12845
rect 16772 12773 16778 12807
rect 16812 12773 16818 12807
rect 16772 12735 16818 12773
rect 16772 12701 16778 12735
rect 16812 12701 16818 12735
rect 16772 12663 16818 12701
rect 16772 12629 16778 12663
rect 16812 12629 16818 12663
rect 16772 12591 16818 12629
rect 16772 12557 16778 12591
rect 16812 12557 16818 12591
rect 16772 12519 16818 12557
rect 16772 12485 16778 12519
rect 16812 12485 16818 12519
rect 16772 12447 16818 12485
rect 16772 12413 16778 12447
rect 16812 12413 16818 12447
rect 16772 12375 16818 12413
rect 16772 12341 16778 12375
rect 16812 12341 16818 12375
rect 16772 12303 16818 12341
rect 16772 12269 16778 12303
rect 16812 12269 16818 12303
rect 16772 12231 16818 12269
rect 16772 12197 16778 12231
rect 16812 12197 16818 12231
rect 16772 12159 16818 12197
rect 16772 12125 16778 12159
rect 16812 12125 16818 12159
rect 16772 12087 16818 12125
rect 16772 12053 16778 12087
rect 16812 12053 16818 12087
rect 16772 12015 16818 12053
rect 16772 11981 16778 12015
rect 16812 11981 16818 12015
rect 16772 11943 16818 11981
rect 16772 11909 16778 11943
rect 16812 11909 16818 11943
rect 16772 11871 16818 11909
rect 16772 11837 16778 11871
rect 16812 11837 16818 11871
rect 16772 11799 16818 11837
rect 16772 11765 16778 11799
rect 16812 11765 16818 11799
rect 16772 11727 16818 11765
rect 16772 11693 16778 11727
rect 16812 11693 16818 11727
rect 16772 11655 16818 11693
rect 16772 11621 16778 11655
rect 16812 11621 16818 11655
rect 16772 11583 16818 11621
rect 16772 11549 16778 11583
rect 16812 11549 16818 11583
rect 16772 11511 16818 11549
rect 16772 11477 16778 11511
rect 16812 11477 16818 11511
rect 16772 11439 16818 11477
rect 16772 11405 16778 11439
rect 16812 11405 16818 11439
rect 16772 11367 16818 11405
rect 16772 11333 16778 11367
rect 16812 11333 16818 11367
rect 16772 11295 16818 11333
rect 16772 11261 16778 11295
rect 16812 11261 16818 11295
rect 16772 11223 16818 11261
rect 16772 11189 16778 11223
rect 16812 11189 16818 11223
rect 16772 11151 16818 11189
rect 16772 11117 16778 11151
rect 16812 11117 16818 11151
rect 16772 11101 16818 11117
rect 16771 11070 16818 11101
rect 16860 12951 16906 12956
rect 16860 12917 16866 12951
rect 16900 12917 16906 12951
rect 16860 12879 16906 12917
rect 16860 12845 16866 12879
rect 16900 12845 16906 12879
rect 16860 12807 16906 12845
rect 16860 12773 16866 12807
rect 16900 12773 16906 12807
rect 16860 12735 16906 12773
rect 16860 12701 16866 12735
rect 16900 12701 16906 12735
rect 16860 12663 16906 12701
rect 16860 12629 16866 12663
rect 16900 12629 16906 12663
rect 16860 12591 16906 12629
rect 16860 12557 16866 12591
rect 16900 12557 16906 12591
rect 16860 12519 16906 12557
rect 16860 12485 16866 12519
rect 16900 12485 16906 12519
rect 16860 12447 16906 12485
rect 16860 12413 16866 12447
rect 16900 12413 16906 12447
rect 16860 12375 16906 12413
rect 16860 12341 16866 12375
rect 16900 12341 16906 12375
rect 16860 12303 16906 12341
rect 16860 12269 16866 12303
rect 16900 12269 16906 12303
rect 16860 12231 16906 12269
rect 16860 12197 16866 12231
rect 16900 12197 16906 12231
rect 16860 12159 16906 12197
rect 16860 12125 16866 12159
rect 16900 12125 16906 12159
rect 16860 12087 16906 12125
rect 16860 12053 16866 12087
rect 16900 12053 16906 12087
rect 16860 12015 16906 12053
rect 16860 11981 16866 12015
rect 16900 11981 16906 12015
rect 16860 11943 16906 11981
rect 16860 11909 16866 11943
rect 16900 11909 16906 11943
rect 16860 11871 16906 11909
rect 16860 11837 16866 11871
rect 16900 11837 16906 11871
rect 16860 11799 16906 11837
rect 16860 11765 16866 11799
rect 16900 11765 16906 11799
rect 16860 11727 16906 11765
rect 16860 11693 16866 11727
rect 16900 11693 16906 11727
rect 16860 11655 16906 11693
rect 16860 11621 16866 11655
rect 16900 11621 16906 11655
rect 16860 11583 16906 11621
rect 16860 11549 16866 11583
rect 16900 11549 16906 11583
rect 16860 11511 16906 11549
rect 16860 11477 16866 11511
rect 16900 11477 16906 11511
rect 16860 11439 16906 11477
rect 16860 11405 16866 11439
rect 16900 11405 16906 11439
rect 16860 11367 16906 11405
rect 16860 11333 16866 11367
rect 16900 11333 16906 11367
rect 16860 11295 16906 11333
rect 16860 11261 16866 11295
rect 16900 11261 16906 11295
rect 16860 11223 16906 11261
rect 16860 11189 16866 11223
rect 16900 11189 16906 11223
rect 16860 11151 16906 11189
rect 16860 11117 16866 11151
rect 16900 11117 16906 11151
rect 16860 11070 16906 11117
rect 16948 12951 16994 12989
rect 17030 13036 17092 13066
rect 17030 12984 17035 13036
rect 17087 12984 17092 13036
rect 17030 12954 17092 12984
rect 17124 13049 17176 13070
rect 17212 13065 17258 13070
rect 17124 13023 17170 13049
rect 17124 12989 17130 13023
rect 17164 12989 17170 13023
rect 16948 12917 16954 12951
rect 16988 12917 16994 12951
rect 16948 12879 16994 12917
rect 16948 12845 16954 12879
rect 16988 12845 16994 12879
rect 16948 12807 16994 12845
rect 16948 12773 16954 12807
rect 16988 12773 16994 12807
rect 16948 12735 16994 12773
rect 16948 12701 16954 12735
rect 16988 12701 16994 12735
rect 16948 12663 16994 12701
rect 16948 12629 16954 12663
rect 16988 12629 16994 12663
rect 16948 12591 16994 12629
rect 16948 12557 16954 12591
rect 16988 12557 16994 12591
rect 16948 12519 16994 12557
rect 16948 12485 16954 12519
rect 16988 12485 16994 12519
rect 16948 12447 16994 12485
rect 16948 12413 16954 12447
rect 16988 12413 16994 12447
rect 16948 12375 16994 12413
rect 16948 12341 16954 12375
rect 16988 12341 16994 12375
rect 16948 12303 16994 12341
rect 16948 12269 16954 12303
rect 16988 12269 16994 12303
rect 16948 12231 16994 12269
rect 16948 12197 16954 12231
rect 16988 12197 16994 12231
rect 16948 12159 16994 12197
rect 16948 12125 16954 12159
rect 16988 12125 16994 12159
rect 16948 12087 16994 12125
rect 16948 12053 16954 12087
rect 16988 12053 16994 12087
rect 16948 12015 16994 12053
rect 16948 11981 16954 12015
rect 16988 11981 16994 12015
rect 16948 11943 16994 11981
rect 16948 11909 16954 11943
rect 16988 11909 16994 11943
rect 16948 11871 16994 11909
rect 16948 11837 16954 11871
rect 16988 11837 16994 11871
rect 16948 11799 16994 11837
rect 16948 11765 16954 11799
rect 16988 11765 16994 11799
rect 16948 11727 16994 11765
rect 16948 11693 16954 11727
rect 16988 11693 16994 11727
rect 16948 11655 16994 11693
rect 16948 11621 16954 11655
rect 16988 11621 16994 11655
rect 16948 11583 16994 11621
rect 16948 11549 16954 11583
rect 16988 11549 16994 11583
rect 16948 11511 16994 11549
rect 16948 11477 16954 11511
rect 16988 11477 16994 11511
rect 16948 11439 16994 11477
rect 16948 11405 16954 11439
rect 16988 11405 16994 11439
rect 16948 11367 16994 11405
rect 16948 11333 16954 11367
rect 16988 11333 16994 11367
rect 16948 11295 16994 11333
rect 16948 11261 16954 11295
rect 16988 11261 16994 11295
rect 16948 11223 16994 11261
rect 16948 11189 16954 11223
rect 16988 11189 16994 11223
rect 16948 11151 16994 11189
rect 16948 11117 16954 11151
rect 16988 11117 16994 11151
rect 16771 10970 16817 11070
rect 16596 10924 16817 10970
rect 16948 10971 16994 11117
rect 17036 12951 17082 12954
rect 17036 12917 17042 12951
rect 17076 12917 17082 12951
rect 17036 12879 17082 12917
rect 17036 12845 17042 12879
rect 17076 12845 17082 12879
rect 17036 12807 17082 12845
rect 17036 12773 17042 12807
rect 17076 12773 17082 12807
rect 17036 12735 17082 12773
rect 17036 12701 17042 12735
rect 17076 12701 17082 12735
rect 17036 12663 17082 12701
rect 17036 12629 17042 12663
rect 17076 12629 17082 12663
rect 17036 12591 17082 12629
rect 17036 12557 17042 12591
rect 17076 12557 17082 12591
rect 17036 12519 17082 12557
rect 17036 12485 17042 12519
rect 17076 12485 17082 12519
rect 17036 12447 17082 12485
rect 17036 12413 17042 12447
rect 17076 12413 17082 12447
rect 17036 12375 17082 12413
rect 17036 12341 17042 12375
rect 17076 12341 17082 12375
rect 17036 12303 17082 12341
rect 17036 12269 17042 12303
rect 17076 12269 17082 12303
rect 17036 12231 17082 12269
rect 17036 12197 17042 12231
rect 17076 12197 17082 12231
rect 17036 12159 17082 12197
rect 17036 12125 17042 12159
rect 17076 12125 17082 12159
rect 17036 12087 17082 12125
rect 17036 12053 17042 12087
rect 17076 12053 17082 12087
rect 17036 12015 17082 12053
rect 17036 11981 17042 12015
rect 17076 11981 17082 12015
rect 17036 11943 17082 11981
rect 17036 11909 17042 11943
rect 17076 11909 17082 11943
rect 17036 11871 17082 11909
rect 17036 11837 17042 11871
rect 17076 11837 17082 11871
rect 17036 11799 17082 11837
rect 17036 11765 17042 11799
rect 17076 11765 17082 11799
rect 17036 11727 17082 11765
rect 17036 11693 17042 11727
rect 17076 11693 17082 11727
rect 17036 11655 17082 11693
rect 17036 11621 17042 11655
rect 17076 11621 17082 11655
rect 17036 11583 17082 11621
rect 17036 11549 17042 11583
rect 17076 11549 17082 11583
rect 17036 11511 17082 11549
rect 17036 11477 17042 11511
rect 17076 11477 17082 11511
rect 17036 11439 17082 11477
rect 17036 11405 17042 11439
rect 17076 11405 17082 11439
rect 17036 11367 17082 11405
rect 17036 11333 17042 11367
rect 17076 11333 17082 11367
rect 17036 11295 17082 11333
rect 17036 11261 17042 11295
rect 17076 11261 17082 11295
rect 17036 11223 17082 11261
rect 17036 11189 17042 11223
rect 17076 11189 17082 11223
rect 17036 11151 17082 11189
rect 17036 11117 17042 11151
rect 17076 11117 17082 11151
rect 17036 11070 17082 11117
rect 17124 12951 17170 12989
rect 17204 13033 17269 13065
rect 17204 12981 17211 13033
rect 17263 12981 17269 13033
rect 17204 12951 17269 12981
rect 17300 13040 17351 13070
rect 17300 13023 17346 13040
rect 17300 12989 17306 13023
rect 17340 12989 17346 13023
rect 17300 12951 17346 12989
rect 17381 13038 17446 13070
rect 17381 12986 17388 13038
rect 17440 12986 17446 13038
rect 17381 12956 17446 12986
rect 17476 13023 17522 13070
rect 17476 12989 17482 13023
rect 17516 12989 17522 13023
rect 17124 12917 17130 12951
rect 17164 12917 17170 12951
rect 17124 12879 17170 12917
rect 17124 12845 17130 12879
rect 17164 12845 17170 12879
rect 17124 12807 17170 12845
rect 17124 12773 17130 12807
rect 17164 12773 17170 12807
rect 17124 12735 17170 12773
rect 17124 12701 17130 12735
rect 17164 12701 17170 12735
rect 17124 12663 17170 12701
rect 17124 12629 17130 12663
rect 17164 12629 17170 12663
rect 17124 12591 17170 12629
rect 17124 12557 17130 12591
rect 17164 12557 17170 12591
rect 17124 12519 17170 12557
rect 17124 12485 17130 12519
rect 17164 12485 17170 12519
rect 17124 12447 17170 12485
rect 17124 12413 17130 12447
rect 17164 12413 17170 12447
rect 17124 12375 17170 12413
rect 17124 12341 17130 12375
rect 17164 12341 17170 12375
rect 17124 12303 17170 12341
rect 17124 12269 17130 12303
rect 17164 12269 17170 12303
rect 17124 12231 17170 12269
rect 17124 12197 17130 12231
rect 17164 12197 17170 12231
rect 17124 12159 17170 12197
rect 17124 12125 17130 12159
rect 17164 12125 17170 12159
rect 17124 12087 17170 12125
rect 17124 12053 17130 12087
rect 17164 12053 17170 12087
rect 17124 12015 17170 12053
rect 17124 11981 17130 12015
rect 17164 11981 17170 12015
rect 17124 11943 17170 11981
rect 17124 11909 17130 11943
rect 17164 11909 17170 11943
rect 17124 11871 17170 11909
rect 17124 11837 17130 11871
rect 17164 11837 17170 11871
rect 17124 11799 17170 11837
rect 17124 11765 17130 11799
rect 17164 11765 17170 11799
rect 17124 11727 17170 11765
rect 17124 11693 17130 11727
rect 17164 11693 17170 11727
rect 17124 11655 17170 11693
rect 17124 11621 17130 11655
rect 17164 11621 17170 11655
rect 17124 11583 17170 11621
rect 17124 11549 17130 11583
rect 17164 11549 17170 11583
rect 17124 11511 17170 11549
rect 17124 11477 17130 11511
rect 17164 11477 17170 11511
rect 17124 11439 17170 11477
rect 17124 11405 17130 11439
rect 17164 11405 17170 11439
rect 17124 11367 17170 11405
rect 17124 11333 17130 11367
rect 17164 11333 17170 11367
rect 17124 11295 17170 11333
rect 17124 11261 17130 11295
rect 17164 11261 17170 11295
rect 17124 11223 17170 11261
rect 17124 11189 17130 11223
rect 17164 11189 17170 11223
rect 17124 11151 17170 11189
rect 17124 11117 17130 11151
rect 17164 11117 17170 11151
rect 17124 11102 17170 11117
rect 17123 11070 17170 11102
rect 17212 12917 17218 12951
rect 17252 12917 17258 12951
rect 17212 12879 17258 12917
rect 17212 12845 17218 12879
rect 17252 12845 17258 12879
rect 17212 12807 17258 12845
rect 17212 12773 17218 12807
rect 17252 12773 17258 12807
rect 17212 12735 17258 12773
rect 17212 12701 17218 12735
rect 17252 12701 17258 12735
rect 17212 12663 17258 12701
rect 17212 12629 17218 12663
rect 17252 12629 17258 12663
rect 17212 12591 17258 12629
rect 17212 12557 17218 12591
rect 17252 12557 17258 12591
rect 17212 12519 17258 12557
rect 17212 12485 17218 12519
rect 17252 12485 17258 12519
rect 17212 12447 17258 12485
rect 17212 12413 17218 12447
rect 17252 12413 17258 12447
rect 17212 12375 17258 12413
rect 17212 12341 17218 12375
rect 17252 12341 17258 12375
rect 17212 12303 17258 12341
rect 17212 12269 17218 12303
rect 17252 12269 17258 12303
rect 17212 12231 17258 12269
rect 17212 12197 17218 12231
rect 17252 12197 17258 12231
rect 17212 12159 17258 12197
rect 17212 12125 17218 12159
rect 17252 12125 17258 12159
rect 17212 12087 17258 12125
rect 17212 12053 17218 12087
rect 17252 12053 17258 12087
rect 17212 12015 17258 12053
rect 17212 11981 17218 12015
rect 17252 11981 17258 12015
rect 17212 11943 17258 11981
rect 17212 11909 17218 11943
rect 17252 11909 17258 11943
rect 17212 11871 17258 11909
rect 17212 11837 17218 11871
rect 17252 11837 17258 11871
rect 17212 11799 17258 11837
rect 17212 11765 17218 11799
rect 17252 11765 17258 11799
rect 17212 11727 17258 11765
rect 17212 11693 17218 11727
rect 17252 11693 17258 11727
rect 17212 11655 17258 11693
rect 17212 11621 17218 11655
rect 17252 11621 17258 11655
rect 17212 11583 17258 11621
rect 17212 11549 17218 11583
rect 17252 11549 17258 11583
rect 17212 11511 17258 11549
rect 17212 11477 17218 11511
rect 17252 11477 17258 11511
rect 17212 11439 17258 11477
rect 17212 11405 17218 11439
rect 17252 11405 17258 11439
rect 17212 11367 17258 11405
rect 17212 11333 17218 11367
rect 17252 11333 17258 11367
rect 17212 11295 17258 11333
rect 17212 11261 17218 11295
rect 17252 11261 17258 11295
rect 17212 11223 17258 11261
rect 17212 11189 17218 11223
rect 17252 11189 17258 11223
rect 17212 11151 17258 11189
rect 17212 11117 17218 11151
rect 17252 11117 17258 11151
rect 17212 11070 17258 11117
rect 17300 12917 17306 12951
rect 17340 12917 17346 12951
rect 17300 12879 17346 12917
rect 17300 12845 17306 12879
rect 17340 12845 17346 12879
rect 17300 12807 17346 12845
rect 17300 12773 17306 12807
rect 17340 12773 17346 12807
rect 17300 12735 17346 12773
rect 17300 12701 17306 12735
rect 17340 12701 17346 12735
rect 17300 12663 17346 12701
rect 17300 12629 17306 12663
rect 17340 12629 17346 12663
rect 17300 12591 17346 12629
rect 17300 12557 17306 12591
rect 17340 12557 17346 12591
rect 17300 12519 17346 12557
rect 17300 12485 17306 12519
rect 17340 12485 17346 12519
rect 17300 12447 17346 12485
rect 17300 12413 17306 12447
rect 17340 12413 17346 12447
rect 17300 12375 17346 12413
rect 17300 12341 17306 12375
rect 17340 12341 17346 12375
rect 17300 12303 17346 12341
rect 17300 12269 17306 12303
rect 17340 12269 17346 12303
rect 17300 12231 17346 12269
rect 17300 12197 17306 12231
rect 17340 12197 17346 12231
rect 17300 12159 17346 12197
rect 17300 12125 17306 12159
rect 17340 12125 17346 12159
rect 17300 12087 17346 12125
rect 17300 12053 17306 12087
rect 17340 12053 17346 12087
rect 17300 12015 17346 12053
rect 17300 11981 17306 12015
rect 17340 11981 17346 12015
rect 17300 11943 17346 11981
rect 17300 11909 17306 11943
rect 17340 11909 17346 11943
rect 17300 11871 17346 11909
rect 17300 11837 17306 11871
rect 17340 11837 17346 11871
rect 17300 11799 17346 11837
rect 17300 11765 17306 11799
rect 17340 11765 17346 11799
rect 17300 11727 17346 11765
rect 17300 11693 17306 11727
rect 17340 11693 17346 11727
rect 17300 11655 17346 11693
rect 17300 11621 17306 11655
rect 17340 11621 17346 11655
rect 17300 11583 17346 11621
rect 17300 11549 17306 11583
rect 17340 11549 17346 11583
rect 17300 11511 17346 11549
rect 17300 11477 17306 11511
rect 17340 11477 17346 11511
rect 17300 11439 17346 11477
rect 17300 11405 17306 11439
rect 17340 11405 17346 11439
rect 17300 11367 17346 11405
rect 17300 11333 17306 11367
rect 17340 11333 17346 11367
rect 17300 11295 17346 11333
rect 17300 11261 17306 11295
rect 17340 11261 17346 11295
rect 17300 11223 17346 11261
rect 17300 11189 17306 11223
rect 17340 11189 17346 11223
rect 17300 11151 17346 11189
rect 17300 11117 17306 11151
rect 17340 11117 17346 11151
rect 17300 11093 17346 11117
rect 17388 12951 17434 12956
rect 17388 12917 17394 12951
rect 17428 12917 17434 12951
rect 17388 12879 17434 12917
rect 17388 12845 17394 12879
rect 17428 12845 17434 12879
rect 17388 12807 17434 12845
rect 17388 12773 17394 12807
rect 17428 12773 17434 12807
rect 17388 12735 17434 12773
rect 17388 12701 17394 12735
rect 17428 12701 17434 12735
rect 17388 12663 17434 12701
rect 17388 12629 17394 12663
rect 17428 12629 17434 12663
rect 17388 12591 17434 12629
rect 17388 12557 17394 12591
rect 17428 12557 17434 12591
rect 17388 12519 17434 12557
rect 17388 12485 17394 12519
rect 17428 12485 17434 12519
rect 17388 12447 17434 12485
rect 17388 12413 17394 12447
rect 17428 12413 17434 12447
rect 17388 12375 17434 12413
rect 17388 12341 17394 12375
rect 17428 12341 17434 12375
rect 17388 12303 17434 12341
rect 17388 12269 17394 12303
rect 17428 12269 17434 12303
rect 17388 12231 17434 12269
rect 17388 12197 17394 12231
rect 17428 12197 17434 12231
rect 17388 12159 17434 12197
rect 17388 12125 17394 12159
rect 17428 12125 17434 12159
rect 17388 12087 17434 12125
rect 17388 12053 17394 12087
rect 17428 12053 17434 12087
rect 17388 12015 17434 12053
rect 17388 11981 17394 12015
rect 17428 11981 17434 12015
rect 17388 11943 17434 11981
rect 17388 11909 17394 11943
rect 17428 11909 17434 11943
rect 17388 11871 17434 11909
rect 17388 11837 17394 11871
rect 17428 11837 17434 11871
rect 17388 11799 17434 11837
rect 17388 11765 17394 11799
rect 17428 11765 17434 11799
rect 17388 11727 17434 11765
rect 17388 11693 17394 11727
rect 17428 11693 17434 11727
rect 17388 11655 17434 11693
rect 17388 11621 17394 11655
rect 17428 11621 17434 11655
rect 17388 11583 17434 11621
rect 17388 11549 17394 11583
rect 17428 11549 17434 11583
rect 17388 11511 17434 11549
rect 17388 11477 17394 11511
rect 17428 11477 17434 11511
rect 17388 11439 17434 11477
rect 17388 11405 17394 11439
rect 17428 11405 17434 11439
rect 17388 11367 17434 11405
rect 17388 11333 17394 11367
rect 17428 11333 17434 11367
rect 17388 11295 17434 11333
rect 17388 11261 17394 11295
rect 17428 11261 17434 11295
rect 17388 11223 17434 11261
rect 17388 11189 17394 11223
rect 17428 11189 17434 11223
rect 17388 11151 17434 11189
rect 17388 11117 17394 11151
rect 17428 11117 17434 11151
rect 17300 11070 17347 11093
rect 17388 11070 17434 11117
rect 17476 12951 17522 12989
rect 17476 12917 17482 12951
rect 17516 12917 17522 12951
rect 17476 12879 17522 12917
rect 17476 12845 17482 12879
rect 17516 12845 17522 12879
rect 17476 12807 17522 12845
rect 17476 12773 17482 12807
rect 17516 12773 17522 12807
rect 17476 12735 17522 12773
rect 17476 12701 17482 12735
rect 17516 12701 17522 12735
rect 17476 12663 17522 12701
rect 17476 12629 17482 12663
rect 17516 12629 17522 12663
rect 17476 12591 17522 12629
rect 17476 12557 17482 12591
rect 17516 12557 17522 12591
rect 17476 12519 17522 12557
rect 17476 12485 17482 12519
rect 17516 12485 17522 12519
rect 17476 12447 17522 12485
rect 17476 12413 17482 12447
rect 17516 12413 17522 12447
rect 17476 12375 17522 12413
rect 17476 12341 17482 12375
rect 17516 12341 17522 12375
rect 17476 12303 17522 12341
rect 17476 12269 17482 12303
rect 17516 12269 17522 12303
rect 17476 12231 17522 12269
rect 17476 12197 17482 12231
rect 17516 12197 17522 12231
rect 17476 12159 17522 12197
rect 17476 12125 17482 12159
rect 17516 12125 17522 12159
rect 17476 12087 17522 12125
rect 17476 12053 17482 12087
rect 17516 12053 17522 12087
rect 17476 12015 17522 12053
rect 17476 11981 17482 12015
rect 17516 11981 17522 12015
rect 17476 11943 17522 11981
rect 17476 11909 17482 11943
rect 17516 11909 17522 11943
rect 17476 11871 17522 11909
rect 17476 11837 17482 11871
rect 17516 11837 17522 11871
rect 17476 11799 17522 11837
rect 17476 11765 17482 11799
rect 17516 11765 17522 11799
rect 17476 11727 17522 11765
rect 17476 11693 17482 11727
rect 17516 11693 17522 11727
rect 17476 11655 17522 11693
rect 17476 11621 17482 11655
rect 17516 11621 17522 11655
rect 17476 11583 17522 11621
rect 17476 11549 17482 11583
rect 17516 11549 17522 11583
rect 17476 11511 17522 11549
rect 17476 11477 17482 11511
rect 17516 11477 17522 11511
rect 17476 11439 17522 11477
rect 17476 11405 17482 11439
rect 17516 11405 17522 11439
rect 17476 11367 17522 11405
rect 17476 11333 17482 11367
rect 17516 11333 17522 11367
rect 17476 11295 17522 11333
rect 17476 11261 17482 11295
rect 17516 11261 17522 11295
rect 17476 11223 17522 11261
rect 17476 11189 17482 11223
rect 17516 11189 17522 11223
rect 17476 11151 17522 11189
rect 17476 11117 17482 11151
rect 17516 11117 17522 11151
rect 17123 10971 17169 11070
rect 16948 10925 17169 10971
rect 17301 10971 17347 11070
rect 17476 10971 17522 11117
rect 17301 10925 17522 10971
rect 13467 10861 13597 10886
rect 13467 10827 13514 10861
rect 13548 10827 13597 10861
rect 13467 10368 13597 10827
rect 14482 10701 14702 10924
rect 17342 10846 17482 10894
rect 17342 10812 17395 10846
rect 17429 10812 17482 10846
rect 17342 10784 17482 10812
rect 14482 10667 14503 10701
rect 14537 10667 14575 10701
rect 14609 10667 14647 10701
rect 14681 10667 14702 10701
rect 14482 10634 14702 10667
rect 17264 10620 17570 10784
rect 17264 10376 17287 10620
rect 17531 10376 17570 10620
rect 17264 10356 17570 10376
rect 17795 10632 18052 16884
rect 17795 10388 17830 10632
rect 18010 10388 18052 10632
rect 17795 10364 18052 10388
rect 4162 9687 26614 9766
rect 4162 8419 4231 9687
rect 5563 9672 26614 9687
rect 5563 9654 25268 9672
rect 5563 8972 13929 9654
rect 16915 8972 25268 9654
rect 5563 8419 25268 8972
rect 4162 8404 25268 8419
rect 26536 8404 26614 9672
rect 4162 8342 26614 8404
rect 2149 7451 28685 7576
rect 2149 6375 2335 7451
rect 3667 7441 28685 7451
rect 3667 6375 27185 7441
rect 2149 6365 27185 6375
rect 28517 6365 28685 7441
rect 2149 6246 28685 6365
<< via1 >>
rect 2351 27715 3683 28791
rect 27191 27787 28523 28863
rect 4248 25660 5516 26928
rect 25306 25668 26574 26936
rect 16834 24564 16856 24591
rect 16856 24564 16886 24591
rect 16834 24539 16886 24564
rect 16750 23993 16802 24001
rect 16750 23959 16758 23993
rect 16758 23959 16792 23993
rect 16792 23959 16802 23993
rect 16750 23949 16802 23959
rect 13670 23053 13786 23361
rect 15285 23366 15401 23610
rect 16302 23548 16418 23553
rect 16302 23442 16307 23548
rect 16307 23442 16413 23548
rect 16413 23442 16418 23548
rect 16302 23437 16418 23442
rect 14050 23103 14102 23117
rect 14050 23069 14066 23103
rect 14066 23069 14100 23103
rect 14100 23069 14102 23103
rect 14050 23065 14102 23069
rect 14250 23103 14302 23117
rect 14250 23069 14258 23103
rect 14258 23069 14292 23103
rect 14292 23069 14302 23103
rect 14250 23065 14302 23069
rect 14440 23103 14492 23117
rect 14440 23069 14450 23103
rect 14450 23069 14484 23103
rect 14484 23069 14492 23103
rect 14440 23065 14492 23069
rect 14630 23103 14682 23117
rect 14630 23069 14642 23103
rect 14642 23069 14676 23103
rect 14676 23069 14682 23103
rect 14630 23065 14682 23069
rect 12585 17712 12765 17956
rect 13960 21231 14012 21237
rect 13960 21197 13970 21231
rect 13970 21197 14004 21231
rect 14004 21197 14012 21231
rect 13960 21185 14012 21197
rect 14150 21231 14202 21237
rect 14150 21197 14162 21231
rect 14162 21197 14196 21231
rect 14196 21197 14202 21231
rect 14150 21185 14202 21197
rect 14340 21231 14392 21237
rect 14340 21197 14354 21231
rect 14354 21197 14388 21231
rect 14388 21197 14392 21231
rect 14340 21185 14392 21197
rect 14530 21231 14582 21237
rect 14530 21197 14546 21231
rect 14546 21197 14580 21231
rect 14580 21197 14582 21231
rect 14530 21185 14582 21197
rect 14839 23107 14891 23116
rect 14839 23073 14848 23107
rect 14848 23073 14882 23107
rect 14882 23073 14891 23107
rect 14839 23064 14891 23073
rect 15910 23142 15962 23157
rect 15910 23108 15926 23142
rect 15926 23108 15960 23142
rect 15960 23108 15962 23142
rect 15910 23105 15962 23108
rect 14730 21231 14782 21237
rect 14730 21197 14738 21231
rect 14738 21197 14772 21231
rect 14772 21197 14782 21231
rect 14730 21185 14782 21197
rect 15810 21270 15862 21277
rect 15810 21236 15830 21270
rect 15830 21236 15862 21270
rect 15810 21225 15862 21236
rect 16100 23142 16152 23157
rect 16100 23108 16118 23142
rect 16118 23108 16152 23142
rect 16100 23105 16152 23108
rect 16658 22121 16710 22130
rect 16658 22087 16662 22121
rect 16662 22087 16696 22121
rect 16696 22087 16710 22121
rect 16658 22078 16710 22087
rect 16940 23993 16992 24001
rect 16940 23959 16950 23993
rect 16950 23959 16984 23993
rect 16984 23959 16992 23993
rect 16940 23949 16992 23959
rect 16839 22121 16891 22130
rect 16839 22087 16854 22121
rect 16854 22087 16888 22121
rect 16888 22087 16891 22121
rect 16839 22078 16891 22087
rect 17130 23993 17182 24001
rect 17130 23959 17142 23993
rect 17142 23959 17176 23993
rect 17176 23959 17182 23993
rect 17130 23949 17182 23959
rect 17029 22121 17081 22130
rect 17029 22087 17046 22121
rect 17046 22087 17080 22121
rect 17080 22087 17081 22121
rect 17029 22078 17081 22087
rect 17320 23993 17372 24001
rect 17320 23959 17334 23993
rect 17334 23959 17368 23993
rect 17368 23959 17372 23993
rect 17320 23949 17372 23959
rect 17220 22121 17272 22133
rect 17220 22087 17238 22121
rect 17238 22087 17272 22121
rect 17220 22081 17272 22087
rect 17520 23993 17572 24001
rect 17520 23959 17526 23993
rect 17526 23959 17560 23993
rect 17560 23959 17572 23993
rect 17520 23949 17572 23959
rect 17419 22121 17471 22131
rect 17419 22087 17430 22121
rect 17430 22087 17464 22121
rect 17464 22087 17471 22121
rect 17419 22079 17471 22087
rect 17610 22121 17662 22132
rect 17610 22087 17622 22121
rect 17622 22087 17656 22121
rect 17656 22087 17662 22121
rect 17610 22080 17662 22087
rect 16010 21270 16062 21277
rect 16010 21236 16022 21270
rect 16022 21236 16056 21270
rect 16056 21236 16062 21270
rect 16010 21225 16062 21236
rect 16877 20941 16993 21313
rect 14940 20518 14992 20546
rect 15004 20518 15056 20546
rect 14940 20494 14974 20518
rect 14974 20494 14992 20518
rect 15004 20494 15008 20518
rect 15008 20494 15056 20518
rect 15068 20494 15120 20546
rect 15132 20518 15184 20546
rect 15196 20518 15248 20546
rect 15132 20494 15166 20518
rect 15166 20494 15184 20518
rect 15196 20494 15200 20518
rect 15200 20494 15248 20518
rect 15260 20494 15312 20546
rect 15324 20518 15376 20546
rect 15388 20518 15440 20546
rect 15324 20494 15358 20518
rect 15358 20494 15376 20518
rect 15388 20494 15392 20518
rect 15392 20494 15440 20518
rect 14914 20398 14926 20401
rect 14926 20398 14960 20401
rect 14960 20398 14966 20401
rect 14914 20360 14966 20398
rect 14914 20349 14926 20360
rect 14926 20349 14960 20360
rect 14960 20349 14966 20360
rect 14824 19246 14830 19261
rect 14830 19246 14864 19261
rect 14864 19246 14876 19261
rect 14824 19209 14876 19246
rect 15104 20398 15118 20401
rect 15118 20398 15152 20401
rect 15152 20398 15156 20401
rect 15104 20360 15156 20398
rect 15104 20349 15118 20360
rect 15118 20349 15152 20360
rect 15152 20349 15156 20360
rect 15014 19246 15022 19261
rect 15022 19246 15056 19261
rect 15056 19246 15066 19261
rect 15014 19209 15066 19246
rect 15304 20398 15310 20401
rect 15310 20398 15344 20401
rect 15344 20398 15356 20401
rect 15304 20360 15356 20398
rect 15304 20349 15310 20360
rect 15310 20349 15344 20360
rect 15344 20349 15356 20360
rect 15204 19246 15214 19261
rect 15214 19246 15248 19261
rect 15248 19246 15256 19261
rect 15204 19209 15256 19246
rect 15494 20398 15502 20401
rect 15502 20398 15536 20401
rect 15536 20398 15546 20401
rect 15494 20360 15546 20398
rect 15494 20349 15502 20360
rect 15502 20349 15536 20360
rect 15536 20349 15546 20360
rect 15394 19246 15406 19261
rect 15406 19246 15440 19261
rect 15440 19246 15446 19261
rect 15394 19209 15446 19246
rect 16074 19903 16086 19921
rect 16086 19903 16120 19921
rect 16120 19903 16126 19921
rect 16074 19869 16126 19903
rect 15974 19217 16026 19251
rect 15974 19199 15990 19217
rect 15990 19199 16024 19217
rect 16024 19199 16026 19217
rect 16264 19903 16278 19921
rect 16278 19903 16312 19921
rect 16312 19903 16316 19921
rect 16264 19869 16316 19903
rect 16174 19217 16226 19251
rect 16174 19199 16182 19217
rect 16182 19199 16216 19217
rect 16216 19199 16226 19217
rect 17067 19232 17119 19241
rect 17067 19198 17072 19232
rect 17072 19198 17106 19232
rect 17106 19198 17119 19232
rect 17067 19189 17119 19198
rect 17131 19232 17183 19241
rect 17131 19198 17144 19232
rect 17144 19198 17178 19232
rect 17178 19198 17183 19232
rect 17131 19189 17183 19198
rect 16524 19049 16576 19101
rect 14163 16576 14279 16692
rect 14669 17800 14694 17809
rect 14694 17800 14721 17809
rect 14669 17762 14721 17800
rect 14669 17757 14694 17762
rect 14694 17757 14721 17762
rect 14669 17728 14694 17745
rect 14694 17728 14721 17745
rect 14669 17693 14721 17728
rect 14669 17656 14694 17681
rect 14694 17656 14721 17681
rect 14669 17629 14721 17656
rect 13534 16310 13586 16362
rect 15119 17803 15171 17810
rect 15119 17769 15138 17803
rect 15138 17769 15171 17803
rect 15119 17758 15171 17769
rect 15119 17731 15171 17746
rect 15119 17697 15138 17731
rect 15138 17697 15171 17731
rect 15119 17694 15171 17697
rect 15119 17659 15171 17682
rect 15119 17630 15138 17659
rect 15138 17630 15171 17659
rect 16804 17964 16856 18016
rect 17372 17919 17488 18012
rect 17372 17885 17414 17919
rect 17414 17885 17448 17919
rect 17448 17885 17488 17919
rect 17372 17847 17488 17885
rect 17372 17813 17414 17847
rect 17414 17813 17448 17847
rect 17448 17813 17488 17847
rect 17372 17775 17488 17813
rect 17372 17768 17414 17775
rect 17414 17768 17448 17775
rect 17448 17768 17488 17775
rect 16765 17325 16945 17505
rect 15459 16635 15511 16687
rect 15459 16571 15511 16623
rect 15045 16422 15097 16474
rect 15045 16358 15097 16410
rect 15045 16294 15097 16346
rect 14766 15976 14818 16000
rect 14766 15948 14792 15976
rect 14792 15948 14818 15976
rect 14502 15857 14554 15870
rect 14502 15823 14518 15857
rect 14518 15823 14552 15857
rect 14552 15823 14554 15857
rect 14502 15818 14554 15823
rect 13528 15421 13580 15437
rect 13528 15387 13572 15421
rect 13572 15387 13580 15421
rect 13528 15385 13580 15387
rect 13528 15349 13580 15373
rect 13528 15321 13572 15349
rect 13572 15321 13580 15349
rect 14422 13985 14474 14000
rect 14422 13951 14456 13985
rect 14456 13951 14474 13985
rect 14422 13948 14474 13951
rect 14702 15857 14754 15870
rect 14702 15823 14710 15857
rect 14710 15823 14744 15857
rect 14744 15823 14754 15857
rect 14702 15818 14754 15823
rect 14602 13985 14654 14000
rect 14602 13951 14614 13985
rect 14614 13951 14648 13985
rect 14648 13951 14654 13985
rect 14602 13948 14654 13951
rect 14892 15857 14944 15870
rect 14892 15823 14902 15857
rect 14902 15823 14936 15857
rect 14936 15823 14944 15857
rect 14892 15818 14944 15823
rect 14792 13985 14844 14000
rect 14792 13951 14806 13985
rect 14806 13951 14840 13985
rect 14840 13951 14844 13985
rect 14792 13948 14844 13951
rect 15082 15857 15134 15870
rect 15082 15823 15094 15857
rect 15094 15823 15128 15857
rect 15128 15823 15134 15857
rect 15082 15818 15134 15823
rect 14982 13985 15034 14000
rect 14982 13951 14998 13985
rect 14998 13951 15032 13985
rect 15032 13951 15034 13985
rect 14982 13948 15034 13951
rect 17182 15896 17234 15910
rect 17182 15862 17188 15896
rect 17188 15862 17222 15896
rect 17222 15862 17234 15896
rect 17182 15858 17234 15862
rect 17372 15896 17424 15910
rect 17372 15862 17380 15896
rect 17380 15862 17414 15896
rect 17414 15862 17424 15896
rect 17372 15858 17424 15862
rect 15172 13985 15224 14000
rect 15172 13951 15190 13985
rect 15190 13951 15224 13985
rect 15172 13948 15224 13951
rect 17082 14024 17134 14030
rect 17082 13990 17092 14024
rect 17092 13990 17126 14024
rect 17126 13990 17134 14024
rect 17082 13978 17134 13990
rect 17282 14024 17334 14030
rect 17282 13990 17284 14024
rect 17284 13990 17318 14024
rect 17318 13990 17334 14024
rect 17282 13978 17334 13990
rect 13611 13832 13616 13859
rect 13616 13832 13650 13859
rect 13650 13832 13663 13859
rect 13611 13807 13663 13832
rect 13513 13023 13565 13032
rect 13513 12989 13522 13023
rect 13522 12989 13556 13023
rect 13556 12989 13565 13023
rect 13513 12980 13565 12989
rect 13685 13023 13737 13036
rect 13685 12989 13698 13023
rect 13698 12989 13732 13023
rect 13732 12989 13737 13023
rect 13685 12984 13737 12989
rect 13861 13023 13913 13032
rect 13861 12989 13874 13023
rect 13874 12989 13908 13023
rect 13908 12989 13913 13023
rect 13861 12980 13913 12989
rect 14042 13023 14094 13038
rect 14042 12989 14050 13023
rect 14050 12989 14084 13023
rect 14084 12989 14094 13023
rect 14042 12986 14094 12989
rect 14217 13023 14269 13038
rect 14217 12989 14226 13023
rect 14226 12989 14260 13023
rect 14260 12989 14269 13023
rect 14217 12986 14269 12989
rect 14395 13023 14447 13038
rect 14395 12989 14402 13023
rect 14402 12989 14436 13023
rect 14436 12989 14447 13023
rect 14395 12986 14447 12989
rect 14567 13023 14619 13036
rect 14567 12989 14578 13023
rect 14578 12989 14612 13023
rect 14612 12989 14619 13023
rect 14567 12984 14619 12989
rect 14747 13023 14799 13039
rect 14747 12989 14754 13023
rect 14754 12989 14788 13023
rect 14788 12989 14799 13023
rect 14747 12987 14799 12989
rect 14921 13023 14973 13036
rect 14921 12989 14930 13023
rect 14930 12989 14964 13023
rect 14964 12989 14973 13023
rect 14921 12984 14973 12989
rect 15098 13023 15150 13038
rect 15098 12989 15106 13023
rect 15106 12989 15140 13023
rect 15140 12989 15150 13023
rect 15098 12986 15150 12989
rect 15275 13023 15327 13038
rect 15275 12989 15282 13023
rect 15282 12989 15316 13023
rect 15316 12989 15327 13023
rect 15275 12986 15327 12989
rect 15450 13023 15502 13033
rect 15450 12989 15458 13023
rect 15458 12989 15492 13023
rect 15492 12989 15502 13023
rect 15450 12981 15502 12989
rect 15627 13023 15679 13038
rect 15627 12989 15634 13023
rect 15634 12989 15668 13023
rect 15668 12989 15679 13023
rect 15627 12986 15679 12989
rect 15803 13023 15855 13033
rect 15803 12989 15810 13023
rect 15810 12989 15844 13023
rect 15844 12989 15855 13023
rect 15803 12981 15855 12989
rect 15977 13023 16029 13034
rect 15977 12989 15986 13023
rect 15986 12989 16020 13023
rect 16020 12989 16029 13023
rect 15977 12982 16029 12989
rect 16155 13023 16207 13033
rect 16155 12989 16162 13023
rect 16162 12989 16196 13023
rect 16196 12989 16207 13023
rect 16155 12981 16207 12989
rect 16331 13023 16383 13034
rect 16331 12989 16338 13023
rect 16338 12989 16372 13023
rect 16372 12989 16383 13023
rect 16331 12982 16383 12989
rect 16509 13023 16561 13032
rect 16509 12989 16514 13023
rect 16514 12989 16548 13023
rect 16548 12989 16561 13023
rect 16509 12980 16561 12989
rect 16681 13023 16733 13036
rect 16681 12989 16690 13023
rect 16690 12989 16724 13023
rect 16724 12989 16733 13023
rect 16681 12984 16733 12989
rect 16858 13023 16910 13038
rect 16858 12989 16866 13023
rect 16866 12989 16900 13023
rect 16900 12989 16910 13023
rect 16858 12986 16910 12989
rect 17035 13023 17087 13036
rect 17035 12989 17042 13023
rect 17042 12989 17076 13023
rect 17076 12989 17087 13023
rect 17035 12984 17087 12989
rect 17211 13023 17263 13033
rect 17211 12989 17218 13023
rect 17218 12989 17252 13023
rect 17252 12989 17263 13023
rect 17211 12981 17263 12989
rect 17388 13023 17440 13038
rect 17388 12989 17394 13023
rect 17394 12989 17428 13023
rect 17428 12989 17440 13023
rect 17388 12986 17440 12989
rect 17287 10376 17531 10620
rect 17830 10388 18010 10632
rect 4231 8419 5563 9687
rect 25268 8404 26536 9672
rect 2335 6375 3667 7451
rect 27185 6365 28517 7441
<< metal2 >>
rect 2168 28791 3820 28952
rect 2168 27715 2351 28791
rect 3683 27715 3820 28791
rect 2168 7451 3820 27715
rect 27052 28863 28704 28952
rect 27052 27787 27191 28863
rect 28523 27787 28704 28863
rect 4162 26928 5612 26992
rect 4162 25660 4248 26928
rect 5516 25660 5612 26928
rect 4162 9687 5612 25660
rect 25230 26936 26614 27010
rect 25230 25668 25306 26936
rect 26574 25668 26614 26936
rect 17828 25329 18030 25342
rect 12324 25277 12582 25328
rect 12324 24901 12344 25277
rect 12560 24901 12582 25277
rect 12324 23390 12582 24901
rect 17828 25113 17864 25329
rect 18000 25113 18030 25329
rect 16810 24591 16910 24620
rect 16810 24539 16834 24591
rect 16886 24539 16910 24591
rect 16810 24426 16910 24539
rect 17828 24426 18030 25113
rect 16810 24250 18030 24426
rect 16810 24050 16910 24250
rect 17828 24248 18030 24250
rect 18170 25271 18480 25326
rect 18170 25055 18216 25271
rect 18432 25055 18480 25271
rect 16810 24041 16950 24050
rect 16743 24040 17003 24041
rect 17123 24040 17193 24041
rect 17313 24040 17383 24041
rect 17513 24040 17583 24041
rect 16740 24001 17583 24040
rect 16740 23949 16750 24001
rect 16802 23949 16940 24001
rect 16992 23949 17130 24001
rect 17182 23949 17320 24001
rect 17372 23949 17520 24001
rect 17572 23949 17583 24001
rect 16740 23911 17583 23949
rect 16740 23910 17570 23911
rect 15260 23610 15432 23632
rect 15260 23596 15285 23610
rect 15401 23596 15432 23610
rect 12324 23388 13786 23390
rect 12324 23361 13802 23388
rect 12324 23053 13670 23361
rect 13786 23053 13802 23361
rect 15260 23380 15275 23596
rect 15411 23380 15432 23596
rect 16270 23553 16450 23580
rect 16270 23437 16302 23553
rect 16418 23437 16450 23553
rect 16270 23410 16450 23437
rect 15260 23366 15285 23380
rect 15401 23366 15432 23380
rect 15260 23312 15432 23366
rect 15901 23190 15971 23191
rect 16091 23190 16161 23191
rect 15901 23157 16161 23190
rect 12324 23032 13802 23053
rect 12334 23030 13802 23032
rect 14041 23150 14111 23151
rect 14241 23150 14311 23151
rect 14431 23150 14501 23151
rect 14621 23150 14691 23151
rect 14041 23117 14910 23150
rect 14041 23065 14050 23117
rect 14102 23065 14250 23117
rect 14302 23065 14440 23117
rect 14492 23065 14630 23117
rect 14682 23116 14910 23117
rect 14682 23065 14839 23116
rect 14041 23064 14839 23065
rect 14891 23064 14910 23116
rect 15901 23105 15910 23157
rect 15962 23105 16100 23157
rect 16152 23105 16161 23157
rect 15901 23071 16161 23105
rect 15920 23070 16160 23071
rect 14041 23031 14910 23064
rect 14060 23030 14910 23031
rect 13648 23028 13802 23030
rect 16316 22170 16444 23410
rect 17213 22170 17283 22173
rect 17412 22170 17482 22171
rect 17603 22170 17673 22172
rect 16316 22133 17673 22170
rect 16316 22130 17220 22133
rect 16316 22078 16658 22130
rect 16710 22078 16839 22130
rect 16891 22078 17029 22130
rect 17081 22081 17220 22130
rect 17272 22132 17673 22133
rect 17272 22131 17610 22132
rect 17272 22081 17419 22131
rect 17081 22079 17419 22081
rect 17471 22080 17610 22131
rect 17662 22080 17673 22132
rect 17471 22079 17673 22080
rect 17081 22078 17673 22079
rect 16316 22042 17673 22078
rect 16650 22040 17660 22042
rect 18170 21356 18480 25055
rect 16840 21313 18481 21356
rect 15801 21310 15871 21311
rect 16001 21310 16071 21311
rect 15801 21277 16071 21310
rect 15801 21274 15810 21277
rect 13964 21271 15810 21274
rect 13951 21237 15810 21271
rect 13951 21185 13960 21237
rect 14012 21185 14150 21237
rect 14202 21185 14340 21237
rect 14392 21185 14530 21237
rect 14582 21185 14730 21237
rect 14782 21225 15810 21237
rect 15862 21225 16010 21277
rect 16062 21274 16071 21277
rect 16062 21225 16074 21274
rect 14782 21185 16074 21225
rect 12358 21092 12859 21158
rect 13951 21151 16074 21185
rect 13964 21146 16074 21151
rect 12358 20476 12425 21092
rect 12801 20903 12859 21092
rect 15615 20903 15745 21146
rect 16840 20941 16877 21313
rect 16993 20941 18481 21313
rect 12801 20731 15766 20903
rect 16840 20902 18481 20941
rect 12801 20476 12859 20731
rect 12358 20416 12859 20476
rect 14540 20546 15490 20570
rect 14540 20494 14940 20546
rect 14992 20494 15004 20546
rect 15056 20494 15068 20546
rect 15120 20494 15132 20546
rect 15184 20494 15196 20546
rect 15248 20494 15260 20546
rect 15312 20494 15324 20546
rect 15376 20494 15388 20546
rect 15440 20494 15490 20546
rect 14540 20470 15490 20494
rect 14550 20020 14650 20470
rect 15615 20440 15745 20731
rect 14900 20401 15745 20440
rect 14900 20349 14914 20401
rect 14966 20349 15104 20401
rect 15156 20349 15304 20401
rect 15356 20349 15494 20401
rect 15546 20349 15745 20401
rect 14900 20310 15745 20349
rect 13010 19920 14650 20020
rect 15615 19965 15745 20310
rect 15615 19960 16175 19965
rect 15615 19921 16330 19960
rect 12531 17956 12811 17995
rect 12531 17942 12585 17956
rect 12765 17942 12811 17956
rect 12531 17726 12567 17942
rect 12783 17726 12811 17942
rect 12531 17712 12585 17726
rect 12765 17712 12811 17726
rect 12531 17677 12811 17712
rect 12640 17088 12940 17130
rect 12640 16872 12677 17088
rect 12893 17080 12940 17088
rect 13010 17080 13110 19920
rect 15615 19869 16074 19921
rect 16126 19869 16264 19921
rect 16316 19869 16330 19921
rect 15615 19840 16330 19869
rect 15615 19835 16175 19840
rect 16060 19830 16140 19835
rect 16250 19830 16330 19840
rect 14810 19261 15460 19300
rect 14810 19209 14824 19261
rect 14876 19209 15014 19261
rect 15066 19209 15204 19261
rect 15256 19209 15394 19261
rect 15446 19209 15460 19261
rect 14810 19170 15460 19209
rect 15960 19280 16040 19290
rect 16160 19280 16240 19290
rect 15960 19251 17230 19280
rect 15960 19199 15974 19251
rect 16026 19199 16174 19251
rect 16226 19241 17230 19251
rect 16226 19199 17067 19241
rect 15960 19189 17067 19199
rect 17119 19189 17131 19241
rect 17183 19189 17230 19241
rect 15960 19160 17230 19189
rect 16490 19101 16620 19130
rect 16490 19049 16524 19101
rect 16576 19049 16620 19101
rect 16490 19020 16620 19049
rect 16500 18050 16620 19020
rect 18200 19068 18590 19110
rect 18200 18985 18247 19068
rect 17725 18695 18247 18985
rect 17330 18050 17530 18060
rect 16500 18038 17530 18050
rect 16500 18016 17362 18038
rect 16500 17964 16804 18016
rect 16856 17964 17362 18016
rect 16500 17930 17362 17964
rect 14642 17810 15187 17851
rect 14642 17809 15119 17810
rect 14642 17757 14669 17809
rect 14721 17758 15119 17809
rect 15171 17758 15187 17810
rect 14721 17757 15187 17758
rect 14642 17746 15187 17757
rect 14642 17745 15119 17746
rect 14642 17693 14669 17745
rect 14721 17694 15119 17745
rect 15171 17694 15187 17746
rect 17330 17742 17362 17930
rect 17498 17742 17530 18038
rect 17330 17720 17530 17742
rect 14721 17693 15187 17694
rect 14642 17682 15187 17693
rect 14642 17681 15119 17682
rect 14642 17629 14669 17681
rect 14721 17630 15119 17681
rect 15171 17630 15187 17682
rect 14721 17629 15187 17630
rect 14642 17594 15187 17629
rect 17725 17570 18015 18695
rect 18200 18612 18247 18695
rect 18543 18985 18590 19068
rect 18543 18695 18635 18985
rect 18543 18612 18590 18695
rect 18200 18580 18590 18612
rect 16720 17566 17230 17570
rect 17270 17566 18020 17570
rect 16720 17505 18020 17566
rect 16720 17325 16765 17505
rect 16945 17325 18020 17505
rect 16720 17286 18020 17325
rect 16720 17280 17230 17286
rect 17270 17280 18020 17286
rect 18110 17253 18521 17306
rect 18110 17205 18170 17253
rect 12893 16980 13110 17080
rect 16741 17045 18170 17205
rect 12893 16872 12940 16980
rect 12640 16830 12940 16872
rect 16741 16714 16901 17045
rect 18110 17037 18170 17045
rect 18466 17037 18521 17253
rect 18110 16980 18521 17037
rect 12860 16692 16901 16714
rect 12860 16576 14163 16692
rect 14279 16687 16901 16692
rect 14279 16635 15459 16687
rect 15511 16635 16901 16687
rect 14279 16623 16901 16635
rect 14279 16576 15459 16623
rect 12860 16571 15459 16576
rect 15511 16571 16901 16623
rect 12860 16554 16901 16571
rect 12490 16098 12770 16140
rect 12490 15802 12522 16098
rect 12738 16000 12770 16098
rect 12860 16000 13020 16554
rect 13506 16364 13602 16397
rect 13506 16308 13532 16364
rect 13588 16308 13602 16364
rect 13506 16279 13602 16308
rect 14486 16264 14646 16554
rect 15016 16474 15126 16494
rect 15016 16452 15045 16474
rect 15097 16452 15126 16474
rect 15016 16396 15043 16452
rect 15099 16396 15126 16452
rect 15016 16372 15045 16396
rect 15097 16372 15126 16396
rect 15016 16316 15043 16372
rect 15099 16316 15126 16372
rect 15016 16294 15045 16316
rect 15097 16294 15126 16316
rect 15016 16274 15126 16294
rect 14486 16234 14966 16264
rect 14486 16104 15196 16234
rect 12738 15840 13020 16000
rect 13119 16070 14305 16073
rect 13119 16000 14844 16070
rect 13119 15948 14766 16000
rect 14818 15948 14844 16000
rect 13119 15932 14844 15948
rect 13119 15851 14305 15932
rect 15036 15904 15196 16104
rect 14486 15870 15196 15904
rect 12738 15802 12770 15840
rect 12490 15770 12770 15802
rect 12512 14257 12732 14258
rect 13119 14257 13341 15851
rect 14486 15818 14502 15870
rect 14554 15818 14702 15870
rect 14754 15818 14892 15870
rect 14944 15818 15082 15870
rect 15134 15818 15196 15870
rect 17173 15910 17433 15944
rect 17173 15858 17182 15910
rect 17234 15858 17372 15910
rect 17424 15858 17433 15910
rect 17173 15824 17433 15858
rect 14486 15794 15196 15818
rect 14486 15784 14646 15794
rect 14693 15784 14763 15794
rect 14883 15784 14953 15794
rect 15073 15784 15143 15794
rect 13507 15437 13602 15452
rect 13507 15407 13528 15437
rect 13580 15407 13602 15437
rect 13507 15351 13526 15407
rect 13582 15351 13602 15407
rect 13507 15321 13528 15351
rect 13580 15321 13602 15351
rect 13507 15307 13602 15321
rect 12512 14036 13341 14257
rect 12512 10620 12733 14036
rect 13119 14035 13341 14036
rect 14413 14029 14483 14034
rect 14593 14029 14663 14034
rect 14783 14029 14853 14034
rect 14973 14029 15043 14034
rect 15163 14029 15233 14034
rect 14413 14000 15233 14029
rect 14413 13948 14422 14000
rect 14474 13948 14602 14000
rect 14654 13948 14792 14000
rect 14844 13948 14982 14000
rect 15034 13948 15172 14000
rect 15224 13948 15233 14000
rect 14413 13914 15233 13948
rect 17073 14030 17343 14064
rect 17073 13978 17082 14030
rect 17134 13978 17282 14030
rect 17334 13978 17343 14030
rect 17073 13944 17343 13978
rect 14419 13911 15227 13914
rect 12862 13883 13120 13900
rect 12862 13871 13662 13883
rect 12862 13859 13668 13871
rect 12862 13807 13611 13859
rect 13663 13807 13668 13859
rect 12862 13794 13668 13807
rect 12862 13745 13662 13794
rect 12482 10589 12760 10620
rect 12862 10612 13120 13745
rect 14672 13071 14862 13911
rect 17132 13071 17332 13944
rect 13519 13070 17434 13071
rect 13519 13062 17446 13070
rect 13508 13039 17446 13062
rect 13508 13038 14747 13039
rect 13508 13036 14042 13038
rect 13508 13032 13685 13036
rect 13508 12980 13513 13032
rect 13565 12984 13685 13032
rect 13737 13032 14042 13036
rect 13737 12984 13861 13032
rect 13565 12980 13861 12984
rect 13913 12986 14042 13032
rect 14094 12986 14217 13038
rect 14269 12986 14395 13038
rect 14447 13036 14747 13038
rect 14447 12986 14567 13036
rect 13913 12984 14567 12986
rect 14619 12987 14747 13036
rect 14799 13038 17446 13039
rect 14799 13036 15098 13038
rect 14799 12987 14921 13036
rect 14619 12984 14921 12987
rect 14973 12986 15098 13036
rect 15150 12986 15275 13038
rect 15327 13033 15627 13038
rect 15327 12986 15450 13033
rect 14973 12984 15450 12986
rect 13913 12981 15450 12984
rect 15502 12986 15627 13033
rect 15679 13036 16858 13038
rect 15679 13034 16681 13036
rect 15679 13033 15977 13034
rect 15679 12986 15803 13033
rect 15502 12981 15803 12986
rect 15855 12982 15977 13033
rect 16029 13033 16331 13034
rect 16029 12982 16155 13033
rect 15855 12981 16155 12982
rect 16207 12982 16331 13033
rect 16383 13032 16681 13034
rect 16383 12982 16509 13032
rect 16207 12981 16509 12982
rect 13913 12980 16509 12981
rect 16561 12984 16681 13032
rect 16733 12986 16858 13036
rect 16910 13036 17388 13038
rect 16910 12986 17035 13036
rect 16733 12984 17035 12986
rect 17087 13033 17388 13036
rect 17087 12984 17211 13033
rect 16561 12981 17211 12984
rect 17263 12986 17388 13033
rect 17440 12986 17446 13038
rect 17263 12981 17446 12986
rect 16561 12980 17446 12981
rect 13508 12956 17446 12980
rect 13508 12950 13570 12956
rect 13678 12954 13743 12956
rect 13856 12950 13918 12956
rect 14562 12954 14624 12956
rect 14672 12954 14862 12956
rect 14916 12954 14978 12956
rect 15443 12951 15508 12956
rect 15796 12951 15861 12956
rect 15972 12952 16034 12956
rect 16148 12951 16213 12956
rect 16326 12952 16388 12956
rect 16502 12950 16567 12956
rect 16676 12954 16738 12956
rect 17030 12954 17092 12956
rect 17204 12951 17269 12956
rect 17262 10620 17568 10784
rect 12482 10373 12509 10589
rect 12725 10373 12760 10589
rect 12482 10342 12760 10373
rect 12856 10590 13126 10612
rect 12856 10374 12882 10590
rect 13098 10374 13126 10590
rect 12856 10356 13126 10374
rect 17262 10376 17287 10620
rect 17531 10376 17568 10620
rect 17262 10356 17568 10376
rect 17792 10632 18052 10712
rect 17792 10618 17830 10632
rect 18010 10618 18052 10632
rect 17792 10402 17812 10618
rect 18028 10402 18052 10618
rect 17792 10388 17830 10402
rect 18010 10388 18052 10402
rect 17792 10366 18052 10388
rect 12868 10354 13126 10356
rect 4162 8419 4231 9687
rect 5563 8419 5612 9687
rect 4162 8324 5612 8419
rect 25230 9672 26614 25668
rect 25230 8404 25268 9672
rect 26536 8404 26614 9672
rect 25230 8342 26614 8404
rect 2168 6375 2335 7451
rect 3667 6375 3820 7451
rect 2168 6246 3820 6375
rect 27052 7441 28704 27787
rect 27052 6365 27185 7441
rect 28517 6365 28704 7441
rect 27052 6246 28704 6365
<< via2 >>
rect 12344 24901 12560 25277
rect 17864 25113 18000 25329
rect 18216 25055 18432 25271
rect 15275 23380 15285 23596
rect 15285 23380 15401 23596
rect 15401 23380 15411 23596
rect 12425 20476 12801 21092
rect 12567 17726 12585 17942
rect 12585 17726 12765 17942
rect 12765 17726 12783 17942
rect 12677 16872 12893 17088
rect 17362 18012 17498 18038
rect 17362 17768 17372 18012
rect 17372 17768 17488 18012
rect 17488 17768 17498 18012
rect 17362 17742 17498 17768
rect 18247 18612 18543 19068
rect 18170 17037 18466 17253
rect 12522 15802 12738 16098
rect 13532 16362 13588 16364
rect 13532 16310 13534 16362
rect 13534 16310 13586 16362
rect 13586 16310 13588 16362
rect 13532 16308 13588 16310
rect 15043 16422 15045 16452
rect 15045 16422 15097 16452
rect 15097 16422 15099 16452
rect 15043 16410 15099 16422
rect 15043 16396 15045 16410
rect 15045 16396 15097 16410
rect 15097 16396 15099 16410
rect 15043 16358 15045 16372
rect 15045 16358 15097 16372
rect 15097 16358 15099 16372
rect 15043 16346 15099 16358
rect 15043 16316 15045 16346
rect 15045 16316 15097 16346
rect 15097 16316 15099 16346
rect 13526 15385 13528 15407
rect 13528 15385 13580 15407
rect 13580 15385 13582 15407
rect 13526 15373 13582 15385
rect 13526 15351 13528 15373
rect 13528 15351 13580 15373
rect 13580 15351 13582 15373
rect 12509 10373 12725 10589
rect 12882 10374 13098 10590
rect 17301 10390 17517 10606
rect 17812 10402 17830 10618
rect 17830 10402 18010 10618
rect 18010 10402 18028 10618
<< metal3 >>
rect 17830 25329 18030 25342
rect 11908 24682 12188 25328
rect 12322 25277 12584 25328
rect 12322 24901 12344 25277
rect 12560 24901 12584 25277
rect 17830 25113 17864 25329
rect 18000 25113 18030 25329
rect 17830 25096 18030 25113
rect 18168 25271 18478 25326
rect 18168 25055 18216 25271
rect 18432 25055 18478 25271
rect 18168 25006 18478 25055
rect 12322 24852 12584 24901
rect 11908 24402 12448 24682
rect 12168 23630 12448 24402
rect 12168 23596 15432 23630
rect 12168 23380 15275 23596
rect 15411 23380 15432 23596
rect 12168 23350 15432 23380
rect 12358 21096 12859 21158
rect 12358 20472 12421 21096
rect 12805 20472 12859 21096
rect 12358 20416 12859 20472
rect 18200 19068 18590 19110
rect 18200 19032 18247 19068
rect 18543 19032 18590 19068
rect 18200 18648 18243 19032
rect 18547 18648 18590 19032
rect 18200 18612 18247 18648
rect 18543 18612 18590 18648
rect 18200 18580 18590 18612
rect 17330 18038 17530 18060
rect 17330 18002 17362 18038
rect 17498 18002 17530 18038
rect 12531 17946 12811 17995
rect 12531 17722 12563 17946
rect 12787 17722 12811 17946
rect 12531 17677 12811 17722
rect 17330 17778 17358 18002
rect 17502 17778 17530 18002
rect 17330 17742 17362 17778
rect 17498 17742 17530 17778
rect 17330 17720 17530 17742
rect 18110 17257 18521 17306
rect 12640 17092 12940 17130
rect 12640 16868 12673 17092
rect 12897 16868 12940 17092
rect 18110 17033 18166 17257
rect 18470 17033 18521 17257
rect 18110 16980 18521 17033
rect 12640 16830 12940 16868
rect 18316 16571 18586 16614
rect 18316 16499 18339 16571
rect 15015 16452 18339 16499
rect 15015 16396 15043 16452
rect 15099 16396 18339 16452
rect 13507 16364 13602 16396
rect 13507 16308 13532 16364
rect 13588 16308 13602 16364
rect 12490 16102 12770 16140
rect 12490 15798 12518 16102
rect 12742 15798 12770 16102
rect 12490 15770 12770 15798
rect 13507 15407 13602 16308
rect 15015 16372 18339 16396
rect 15015 16316 15043 16372
rect 15099 16316 18339 16372
rect 15015 16288 18339 16316
rect 15016 16274 15126 16288
rect 18316 16267 18339 16288
rect 18563 16267 18586 16571
rect 18316 16224 18586 16267
rect 13507 15351 13526 15407
rect 13582 15351 13602 15407
rect 13507 15307 13602 15351
rect 12482 10589 12760 10620
rect 17262 10606 17568 10784
rect 12482 10373 12509 10589
rect 12725 10373 12760 10589
rect 12482 10342 12760 10373
rect 12862 10590 13120 10604
rect 12862 10374 12882 10590
rect 13098 10374 13120 10590
rect 12862 10360 13120 10374
rect 17262 10390 17301 10606
rect 17517 10390 17568 10606
rect 17262 10356 17568 10390
rect 17792 10618 18052 10712
rect 17792 10402 17812 10618
rect 18028 10402 18052 10618
rect 17792 10366 18052 10402
<< via3 >>
rect 12421 21092 12805 21096
rect 12421 20476 12425 21092
rect 12425 20476 12801 21092
rect 12801 20476 12805 21092
rect 12421 20472 12805 20476
rect 18243 18648 18247 19032
rect 18247 18648 18543 19032
rect 18543 18648 18547 19032
rect 12563 17942 12787 17946
rect 12563 17726 12567 17942
rect 12567 17726 12783 17942
rect 12783 17726 12787 17942
rect 12563 17722 12787 17726
rect 17358 17778 17362 18002
rect 17362 17778 17498 18002
rect 17498 17778 17502 18002
rect 12673 17088 12897 17092
rect 12673 16872 12677 17088
rect 12677 16872 12893 17088
rect 12893 16872 12897 17088
rect 12673 16868 12897 16872
rect 18166 17253 18470 17257
rect 18166 17037 18170 17253
rect 18170 17037 18466 17253
rect 18466 17037 18470 17253
rect 18166 17033 18470 17037
rect 12518 16098 12742 16102
rect 12518 15802 12522 16098
rect 12522 15802 12738 16098
rect 12738 15802 12742 16098
rect 12518 15798 12742 15802
rect 18339 16267 18563 16571
<< metal4 >>
rect 5947 17996 12147 24400
rect 12358 21096 12859 21158
rect 12358 20472 12421 21096
rect 12805 20472 12859 21096
rect 12358 20416 12859 20472
rect 18200 19032 18590 19110
rect 18200 18648 18243 19032
rect 18547 18648 18590 19032
rect 18200 18580 18590 18648
rect 18861 18060 25061 24454
rect 17330 18008 25061 18060
rect 17330 18002 18963 18008
rect 5947 17954 12813 17996
rect 5947 17718 6049 17954
rect 6285 17718 6369 17954
rect 6605 17718 6689 17954
rect 6925 17718 7009 17954
rect 7245 17718 7329 17954
rect 7565 17718 7649 17954
rect 7885 17718 7969 17954
rect 8205 17718 8289 17954
rect 8525 17718 8609 17954
rect 8845 17718 8929 17954
rect 9165 17718 9249 17954
rect 9485 17718 9569 17954
rect 9805 17718 9889 17954
rect 10125 17718 10209 17954
rect 10445 17718 10529 17954
rect 10765 17718 10849 17954
rect 11085 17718 11169 17954
rect 11405 17718 11489 17954
rect 11725 17718 11809 17954
rect 12045 17946 12813 17954
rect 12045 17722 12563 17946
rect 12787 17722 12813 17946
rect 12045 17718 12813 17722
rect 17330 17778 17358 18002
rect 17502 17778 18963 18002
rect 17330 17772 18963 17778
rect 19199 17772 19283 18008
rect 19519 17772 19603 18008
rect 19839 17772 19923 18008
rect 20159 17772 20243 18008
rect 20479 17772 20563 18008
rect 20799 17772 20883 18008
rect 21119 17772 21203 18008
rect 21439 17772 21523 18008
rect 21759 17772 21843 18008
rect 22079 17772 22163 18008
rect 22399 17772 22483 18008
rect 22719 17772 22803 18008
rect 23039 17772 23123 18008
rect 23359 17772 23443 18008
rect 23679 17772 23763 18008
rect 23999 17772 24083 18008
rect 24319 17772 24403 18008
rect 24639 17772 24723 18008
rect 24959 17772 25061 18008
rect 17330 17752 25061 17772
rect 17330 17720 19240 17752
rect 5947 17698 12813 17718
rect 11905 17677 12813 17698
rect 18110 17282 19228 17305
rect 18110 17262 25060 17282
rect 18110 17257 18962 17262
rect 5991 17130 12191 17132
rect 5991 17112 12940 17130
rect 5991 16876 6093 17112
rect 6329 16876 6413 17112
rect 6649 16876 6733 17112
rect 6969 16876 7053 17112
rect 7289 16876 7373 17112
rect 7609 16876 7693 17112
rect 7929 16876 8013 17112
rect 8249 16876 8333 17112
rect 8569 16876 8653 17112
rect 8889 16876 8973 17112
rect 9209 16876 9293 17112
rect 9529 16876 9613 17112
rect 9849 16876 9933 17112
rect 10169 16876 10253 17112
rect 10489 16876 10573 17112
rect 10809 16876 10893 17112
rect 11129 16876 11213 17112
rect 11449 16876 11533 17112
rect 11769 16876 11853 17112
rect 12089 17092 12940 17112
rect 12089 16876 12673 17092
rect 5991 16868 12673 16876
rect 12897 16868 12940 17092
rect 18110 17033 18166 17257
rect 18470 17033 18962 17257
rect 18110 17026 18962 17033
rect 19198 17026 19282 17262
rect 19518 17026 19602 17262
rect 19838 17026 19922 17262
rect 20158 17026 20242 17262
rect 20478 17026 20562 17262
rect 20798 17026 20882 17262
rect 21118 17026 21202 17262
rect 21438 17026 21522 17262
rect 21758 17026 21842 17262
rect 22078 17026 22162 17262
rect 22398 17026 22482 17262
rect 22718 17026 22802 17262
rect 23038 17026 23122 17262
rect 23358 17026 23442 17262
rect 23678 17026 23762 17262
rect 23998 17026 24082 17262
rect 24318 17026 24402 17262
rect 24638 17026 24722 17262
rect 24958 17026 25060 17262
rect 18110 16980 25060 17026
rect 5991 16830 12940 16868
rect 5991 10430 12191 16830
rect 18316 16571 18586 16614
rect 18316 16536 18339 16571
rect 18563 16536 18586 16571
rect 18316 16300 18334 16536
rect 18570 16300 18586 16536
rect 18316 16267 18339 16300
rect 18563 16267 18586 16300
rect 18316 16224 18586 16267
rect 12490 16102 12770 16140
rect 12490 16068 12518 16102
rect 12742 16068 12770 16102
rect 12490 15832 12512 16068
rect 12748 15832 12770 16068
rect 12490 15798 12518 15832
rect 12742 15798 12770 15832
rect 12490 15770 12770 15798
rect 18860 10580 25060 16980
<< via4 >>
rect 12495 20826 12731 21062
rect 12495 20506 12731 20742
rect 18277 18722 18513 18958
rect 6049 17718 6285 17954
rect 6369 17718 6605 17954
rect 6689 17718 6925 17954
rect 7009 17718 7245 17954
rect 7329 17718 7565 17954
rect 7649 17718 7885 17954
rect 7969 17718 8205 17954
rect 8289 17718 8525 17954
rect 8609 17718 8845 17954
rect 8929 17718 9165 17954
rect 9249 17718 9485 17954
rect 9569 17718 9805 17954
rect 9889 17718 10125 17954
rect 10209 17718 10445 17954
rect 10529 17718 10765 17954
rect 10849 17718 11085 17954
rect 11169 17718 11405 17954
rect 11489 17718 11725 17954
rect 11809 17718 12045 17954
rect 18963 17772 19199 18008
rect 19283 17772 19519 18008
rect 19603 17772 19839 18008
rect 19923 17772 20159 18008
rect 20243 17772 20479 18008
rect 20563 17772 20799 18008
rect 20883 17772 21119 18008
rect 21203 17772 21439 18008
rect 21523 17772 21759 18008
rect 21843 17772 22079 18008
rect 22163 17772 22399 18008
rect 22483 17772 22719 18008
rect 22803 17772 23039 18008
rect 23123 17772 23359 18008
rect 23443 17772 23679 18008
rect 23763 17772 23999 18008
rect 24083 17772 24319 18008
rect 24403 17772 24639 18008
rect 24723 17772 24959 18008
rect 6093 16876 6329 17112
rect 6413 16876 6649 17112
rect 6733 16876 6969 17112
rect 7053 16876 7289 17112
rect 7373 16876 7609 17112
rect 7693 16876 7929 17112
rect 8013 16876 8249 17112
rect 8333 16876 8569 17112
rect 8653 16876 8889 17112
rect 8973 16876 9209 17112
rect 9293 16876 9529 17112
rect 9613 16876 9849 17112
rect 9933 16876 10169 17112
rect 10253 16876 10489 17112
rect 10573 16876 10809 17112
rect 10893 16876 11129 17112
rect 11213 16876 11449 17112
rect 11533 16876 11769 17112
rect 11853 16876 12089 17112
rect 18962 17026 19198 17262
rect 19282 17026 19518 17262
rect 19602 17026 19838 17262
rect 19922 17026 20158 17262
rect 20242 17026 20478 17262
rect 20562 17026 20798 17262
rect 20882 17026 21118 17262
rect 21202 17026 21438 17262
rect 21522 17026 21758 17262
rect 21842 17026 22078 17262
rect 22162 17026 22398 17262
rect 22482 17026 22718 17262
rect 22802 17026 23038 17262
rect 23122 17026 23358 17262
rect 23442 17026 23678 17262
rect 23762 17026 23998 17262
rect 24082 17026 24318 17262
rect 24402 17026 24638 17262
rect 24722 17026 24958 17262
rect 18334 16300 18339 16536
rect 18339 16300 18563 16536
rect 18563 16300 18570 16536
rect 12512 15832 12518 16068
rect 12518 15832 12742 16068
rect 12742 15832 12748 16068
<< mimcap2 >>
rect 6047 24138 12047 24300
rect 6047 18462 6209 24138
rect 11885 18462 12047 24138
rect 6047 18300 12047 18462
rect 18961 24192 24961 24354
rect 18961 18516 19123 24192
rect 24799 18516 24961 24192
rect 18961 18354 24961 18516
rect 6091 16368 12091 16530
rect 6091 10692 6253 16368
rect 11929 10692 12091 16368
rect 6091 10530 12091 10692
rect 18960 16518 24960 16680
rect 18960 10842 19122 16518
rect 24798 10842 24960 16518
rect 18960 10680 24960 10842
<< mimcap2contact >>
rect 6209 18462 11885 24138
rect 19123 18516 24799 24192
rect 6253 10692 11929 16368
rect 19122 10842 24798 16518
<< metal5 >>
rect 6063 24138 12031 24284
rect 6063 18462 6209 24138
rect 11885 21154 12031 24138
rect 18977 24192 24945 24338
rect 11885 21062 12857 21154
rect 11885 20826 12495 21062
rect 12731 20826 12857 21062
rect 11885 20742 12857 20826
rect 11885 20506 12495 20742
rect 12731 20506 12857 20742
rect 11885 20418 12857 20506
rect 11885 18462 12031 20418
rect 18977 19110 19123 24192
rect 18200 18958 19123 19110
rect 18200 18722 18277 18958
rect 18513 18722 19123 18958
rect 18200 18580 19123 18722
rect 6063 18316 12031 18462
rect 18977 18516 19123 18580
rect 24799 18516 24945 24192
rect 18977 18370 24945 18516
rect 18860 18008 25062 18050
rect 5946 17954 12148 17996
rect 5946 17718 6049 17954
rect 6285 17718 6369 17954
rect 6605 17718 6689 17954
rect 6925 17718 7009 17954
rect 7245 17718 7329 17954
rect 7565 17718 7649 17954
rect 7885 17718 7969 17954
rect 8205 17718 8289 17954
rect 8525 17718 8609 17954
rect 8845 17718 8929 17954
rect 9165 17718 9249 17954
rect 9485 17718 9569 17954
rect 9805 17718 9889 17954
rect 10125 17718 10209 17954
rect 10445 17718 10529 17954
rect 10765 17718 10849 17954
rect 11085 17718 11169 17954
rect 11405 17718 11489 17954
rect 11725 17718 11809 17954
rect 12045 17718 12148 17954
rect 18860 17772 18963 18008
rect 19199 17772 19283 18008
rect 19519 17772 19603 18008
rect 19839 17772 19923 18008
rect 20159 17772 20243 18008
rect 20479 17772 20563 18008
rect 20799 17772 20883 18008
rect 21119 17772 21203 18008
rect 21439 17772 21523 18008
rect 21759 17772 21843 18008
rect 22079 17772 22163 18008
rect 22399 17772 22483 18008
rect 22719 17772 22803 18008
rect 23039 17772 23123 18008
rect 23359 17772 23443 18008
rect 23679 17772 23763 18008
rect 23999 17772 24083 18008
rect 24319 17772 24403 18008
rect 24639 17772 24723 18008
rect 24959 17772 25062 18008
rect 18860 17730 25062 17772
rect 5946 17676 12148 17718
rect 18859 17262 25061 17304
rect 5990 17112 12192 17154
rect 5990 16876 6093 17112
rect 6329 16876 6413 17112
rect 6649 16876 6733 17112
rect 6969 16876 7053 17112
rect 7289 16876 7373 17112
rect 7609 16876 7693 17112
rect 7929 16876 8013 17112
rect 8249 16876 8333 17112
rect 8569 16876 8653 17112
rect 8889 16876 8973 17112
rect 9209 16876 9293 17112
rect 9529 16876 9613 17112
rect 9849 16876 9933 17112
rect 10169 16876 10253 17112
rect 10489 16876 10573 17112
rect 10809 16876 10893 17112
rect 11129 16876 11213 17112
rect 11449 16876 11533 17112
rect 11769 16876 11853 17112
rect 12089 16876 12192 17112
rect 18859 17026 18962 17262
rect 19198 17026 19282 17262
rect 19518 17026 19602 17262
rect 19838 17026 19922 17262
rect 20158 17026 20242 17262
rect 20478 17026 20562 17262
rect 20798 17026 20882 17262
rect 21118 17026 21202 17262
rect 21438 17026 21522 17262
rect 21758 17026 21842 17262
rect 22078 17026 22162 17262
rect 22398 17026 22482 17262
rect 22718 17026 22802 17262
rect 23038 17026 23122 17262
rect 23358 17026 23442 17262
rect 23678 17026 23762 17262
rect 23998 17026 24082 17262
rect 24318 17026 24402 17262
rect 24638 17026 24722 17262
rect 24958 17026 25061 17262
rect 18859 16984 25061 17026
rect 5990 16834 12192 16876
rect 18976 16614 24944 16664
rect 18281 16536 24944 16614
rect 6107 16368 12075 16514
rect 6107 10692 6253 16368
rect 11929 16160 12075 16368
rect 18281 16300 18334 16536
rect 18570 16518 24944 16536
rect 18570 16300 19122 16518
rect 18281 16224 19122 16300
rect 11929 16068 12800 16160
rect 11929 15832 12512 16068
rect 12748 15832 12800 16068
rect 11929 15750 12800 15832
rect 11929 10692 12075 15750
rect 18976 10842 19122 16224
rect 24798 10842 24944 16518
rect 18976 10696 24944 10842
rect 6107 10546 12075 10692
<< labels >>
flabel metal1 s 13514 10494 13514 10494 0 FreeSans 2000 90 0 0 VRF
port 1 nsew
flabel locali s 15294 10468 15294 10468 0 FreeSans 1600 90 0 0 VSS
port 2 nsew
flabel metal3 s 13002 10468 13002 10468 0 FreeSans 1600 90 0 0 VB0_75
port 3 nsew
flabel metal3 s 17420 10482 17420 10482 0 FreeSans 1600 90 0 0 VSI1
port 4 nsew
flabel metal3 s 12582 10524 12582 10524 0 FreeSans 1600 90 0 0 VB1_4
port 5 nsew
flabel locali s 14542 25052 14542 25052 0 FreeSans 1600 90 0 0 VDD
port 6 nsew
flabel metal3 s 17906 10532 17906 10532 0 FreeSans 1600 90 0 0 VB1_5
port 7 nsew
flabel metal3 s 18282 25126 18282 25126 0 FreeSans 1600 90 0 0 VB0_9
port 8 nsew
flabel metal3 s 12442 25032 12442 25032 0 FreeSans 1600 90 0 0 VSI2
port 9 nsew
flabel metal3 s 12000 25086 12000 25086 0 FreeSans 1600 90 0 0 VB0_6
port 10 nsew
flabel metal3 s 17928 25256 17928 25256 0 FreeSans 1600 90 0 0 VOUT
port 11 nsew
<< end >>
