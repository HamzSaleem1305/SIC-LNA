magic
tech sky130A
magscale 1 2
timestamp 1666420471
<< pwell >>
rect -201 -998 201 998
<< psubdiff >>
rect -165 928 -69 962
rect 69 928 165 962
rect -165 866 -131 928
rect 131 866 165 928
rect -165 -928 -131 -866
rect 131 -928 165 -866
rect -165 -962 -69 -928
rect 69 -962 165 -928
<< psubdiffcont >>
rect -69 928 69 962
rect -165 -866 -131 866
rect 131 -866 165 866
rect -69 -962 69 -928
<< xpolycontact >>
rect -35 400 35 832
rect -35 -832 35 -400
<< ppolyres >>
rect -35 -400 35 400
<< locali >>
rect -165 928 -69 962
rect 69 928 165 962
rect -165 866 -131 928
rect 131 866 165 928
rect -165 -928 -131 -866
rect 131 -928 165 -866
rect -165 -962 -69 -928
rect 69 -962 165 -928
<< viali >>
rect -19 417 19 814
rect -19 -814 19 -417
<< metal1 >>
rect -25 814 25 826
rect -25 417 -19 814
rect 19 417 25 814
rect -25 405 25 417
rect -25 -417 25 -405
rect -25 -814 -19 -417
rect 19 -814 25 -417
rect -25 -826 25 -814
<< res0p35 >>
rect -37 -402 37 402
<< properties >>
string FIXED_BBOX -148 -945 148 945
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 4 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 3.764k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
