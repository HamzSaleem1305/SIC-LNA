magic
tech sky130A
timestamp 1640952342
<< error_p >>
rect -72 -741 72 741
<< nwell >>
rect -72 -741 72 741
<< pmoslvt >>
rect -25 -710 25 710
<< pdiff >>
rect -54 704 -25 710
rect -54 -704 -48 704
rect -31 -704 -25 704
rect -54 -710 -25 -704
rect 25 704 54 710
rect 25 -704 31 704
rect 48 -704 54 704
rect 25 -710 54 -704
<< pdiffc >>
rect -48 -704 -31 704
rect 31 -704 48 704
<< poly >>
rect -25 710 25 723
rect -25 -723 25 -710
<< locali >>
rect -48 704 -31 712
rect -48 -712 -31 -704
rect 31 704 48 712
rect 31 -712 48 -704
<< viali >>
rect -48 -704 -31 704
rect 31 -704 48 704
<< metal1 >>
rect -51 704 -28 710
rect -51 -704 -48 704
rect -31 -704 -28 704
rect -51 -710 -28 -704
rect 28 704 51 710
rect 28 -704 31 704
rect 48 -704 51 704
rect 28 -710 51 -704
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 14.2 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
