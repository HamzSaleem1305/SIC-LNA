magic
tech sky130A
magscale 1 2
timestamp 1666360620
<< error_p >>
rect -941 1072 -883 1078
rect -749 1072 -691 1078
rect -557 1072 -499 1078
rect -365 1072 -307 1078
rect -173 1072 -115 1078
rect 19 1072 77 1078
rect 211 1072 269 1078
rect 403 1072 461 1078
rect 595 1072 653 1078
rect 787 1072 845 1078
rect 979 1072 1037 1078
rect -941 1038 -929 1072
rect -749 1038 -737 1072
rect -557 1038 -545 1072
rect -365 1038 -353 1072
rect -173 1038 -161 1072
rect 19 1038 31 1072
rect 211 1038 223 1072
rect 403 1038 415 1072
rect 595 1038 607 1072
rect 787 1038 799 1072
rect 979 1038 991 1072
rect -941 1032 -883 1038
rect -749 1032 -691 1038
rect -557 1032 -499 1038
rect -365 1032 -307 1038
rect -173 1032 -115 1038
rect 19 1032 77 1038
rect 211 1032 269 1038
rect 403 1032 461 1038
rect 595 1032 653 1038
rect 787 1032 845 1038
rect 979 1032 1037 1038
rect -1037 -1038 -979 -1032
rect -845 -1038 -787 -1032
rect -653 -1038 -595 -1032
rect -461 -1038 -403 -1032
rect -269 -1038 -211 -1032
rect -77 -1038 -19 -1032
rect 115 -1038 173 -1032
rect 307 -1038 365 -1032
rect 499 -1038 557 -1032
rect 691 -1038 749 -1032
rect 883 -1038 941 -1032
rect -1037 -1072 -1025 -1038
rect -845 -1072 -833 -1038
rect -653 -1072 -641 -1038
rect -461 -1072 -449 -1038
rect -269 -1072 -257 -1038
rect -77 -1072 -65 -1038
rect 115 -1072 127 -1038
rect 307 -1072 319 -1038
rect 499 -1072 511 -1038
rect 691 -1072 703 -1038
rect 883 -1072 895 -1038
rect -1037 -1078 -979 -1072
rect -845 -1078 -787 -1072
rect -653 -1078 -595 -1072
rect -461 -1078 -403 -1072
rect -269 -1078 -211 -1072
rect -77 -1078 -19 -1072
rect 115 -1078 173 -1072
rect 307 -1078 365 -1072
rect 499 -1078 557 -1072
rect 691 -1078 749 -1072
rect 883 -1078 941 -1072
<< pwell >>
rect -1223 -1210 1223 1210
<< nmoslvt >>
rect -1023 -1000 -993 1000
rect -927 -1000 -897 1000
rect -831 -1000 -801 1000
rect -735 -1000 -705 1000
rect -639 -1000 -609 1000
rect -543 -1000 -513 1000
rect -447 -1000 -417 1000
rect -351 -1000 -321 1000
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
rect 321 -1000 351 1000
rect 417 -1000 447 1000
rect 513 -1000 543 1000
rect 609 -1000 639 1000
rect 705 -1000 735 1000
rect 801 -1000 831 1000
rect 897 -1000 927 1000
rect 993 -1000 1023 1000
<< ndiff >>
rect -1085 988 -1023 1000
rect -1085 -988 -1073 988
rect -1039 -988 -1023 988
rect -1085 -1000 -1023 -988
rect -993 988 -927 1000
rect -993 -988 -977 988
rect -943 -988 -927 988
rect -993 -1000 -927 -988
rect -897 988 -831 1000
rect -897 -988 -881 988
rect -847 -988 -831 988
rect -897 -1000 -831 -988
rect -801 988 -735 1000
rect -801 -988 -785 988
rect -751 -988 -735 988
rect -801 -1000 -735 -988
rect -705 988 -639 1000
rect -705 -988 -689 988
rect -655 -988 -639 988
rect -705 -1000 -639 -988
rect -609 988 -543 1000
rect -609 -988 -593 988
rect -559 -988 -543 988
rect -609 -1000 -543 -988
rect -513 988 -447 1000
rect -513 -988 -497 988
rect -463 -988 -447 988
rect -513 -1000 -447 -988
rect -417 988 -351 1000
rect -417 -988 -401 988
rect -367 -988 -351 988
rect -417 -1000 -351 -988
rect -321 988 -255 1000
rect -321 -988 -305 988
rect -271 -988 -255 988
rect -321 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 321 1000
rect 255 -988 271 988
rect 305 -988 321 988
rect 255 -1000 321 -988
rect 351 988 417 1000
rect 351 -988 367 988
rect 401 -988 417 988
rect 351 -1000 417 -988
rect 447 988 513 1000
rect 447 -988 463 988
rect 497 -988 513 988
rect 447 -1000 513 -988
rect 543 988 609 1000
rect 543 -988 559 988
rect 593 -988 609 988
rect 543 -1000 609 -988
rect 639 988 705 1000
rect 639 -988 655 988
rect 689 -988 705 988
rect 639 -1000 705 -988
rect 735 988 801 1000
rect 735 -988 751 988
rect 785 -988 801 988
rect 735 -1000 801 -988
rect 831 988 897 1000
rect 831 -988 847 988
rect 881 -988 897 988
rect 831 -1000 897 -988
rect 927 988 993 1000
rect 927 -988 943 988
rect 977 -988 993 988
rect 927 -1000 993 -988
rect 1023 988 1085 1000
rect 1023 -988 1039 988
rect 1073 -988 1085 988
rect 1023 -1000 1085 -988
<< ndiffc >>
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
<< psubdiff >>
rect -1187 1140 -1091 1174
rect 1091 1140 1187 1174
rect -1187 1078 -1153 1140
rect 1153 1078 1187 1140
rect -1187 -1140 -1153 -1078
rect 1153 -1140 1187 -1078
rect -1187 -1174 -1091 -1140
rect 1091 -1174 1187 -1140
<< psubdiffcont >>
rect -1091 1140 1091 1174
rect -1187 -1078 -1153 1078
rect 1153 -1078 1187 1078
rect -1091 -1174 1091 -1140
<< poly >>
rect -945 1072 -879 1088
rect -945 1038 -929 1072
rect -895 1038 -879 1072
rect -1023 1000 -993 1026
rect -945 1022 -879 1038
rect -753 1072 -687 1088
rect -753 1038 -737 1072
rect -703 1038 -687 1072
rect -927 1000 -897 1022
rect -831 1000 -801 1026
rect -753 1022 -687 1038
rect -561 1072 -495 1088
rect -561 1038 -545 1072
rect -511 1038 -495 1072
rect -735 1000 -705 1022
rect -639 1000 -609 1026
rect -561 1022 -495 1038
rect -369 1072 -303 1088
rect -369 1038 -353 1072
rect -319 1038 -303 1072
rect -543 1000 -513 1022
rect -447 1000 -417 1026
rect -369 1022 -303 1038
rect -177 1072 -111 1088
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect -351 1000 -321 1022
rect -255 1000 -225 1026
rect -177 1022 -111 1038
rect 15 1072 81 1088
rect 15 1038 31 1072
rect 65 1038 81 1072
rect -159 1000 -129 1022
rect -63 1000 -33 1026
rect 15 1022 81 1038
rect 207 1072 273 1088
rect 207 1038 223 1072
rect 257 1038 273 1072
rect 33 1000 63 1022
rect 129 1000 159 1026
rect 207 1022 273 1038
rect 399 1072 465 1088
rect 399 1038 415 1072
rect 449 1038 465 1072
rect 225 1000 255 1022
rect 321 1000 351 1026
rect 399 1022 465 1038
rect 591 1072 657 1088
rect 591 1038 607 1072
rect 641 1038 657 1072
rect 417 1000 447 1022
rect 513 1000 543 1026
rect 591 1022 657 1038
rect 783 1072 849 1088
rect 783 1038 799 1072
rect 833 1038 849 1072
rect 609 1000 639 1022
rect 705 1000 735 1026
rect 783 1022 849 1038
rect 975 1072 1041 1088
rect 975 1038 991 1072
rect 1025 1038 1041 1072
rect 801 1000 831 1022
rect 897 1000 927 1026
rect 975 1022 1041 1038
rect 993 1000 1023 1022
rect -1023 -1022 -993 -1000
rect -1041 -1038 -975 -1022
rect -927 -1026 -897 -1000
rect -831 -1022 -801 -1000
rect -1041 -1072 -1025 -1038
rect -991 -1072 -975 -1038
rect -1041 -1088 -975 -1072
rect -849 -1038 -783 -1022
rect -735 -1026 -705 -1000
rect -639 -1022 -609 -1000
rect -849 -1072 -833 -1038
rect -799 -1072 -783 -1038
rect -849 -1088 -783 -1072
rect -657 -1038 -591 -1022
rect -543 -1026 -513 -1000
rect -447 -1022 -417 -1000
rect -657 -1072 -641 -1038
rect -607 -1072 -591 -1038
rect -657 -1088 -591 -1072
rect -465 -1038 -399 -1022
rect -351 -1026 -321 -1000
rect -255 -1022 -225 -1000
rect -465 -1072 -449 -1038
rect -415 -1072 -399 -1038
rect -465 -1088 -399 -1072
rect -273 -1038 -207 -1022
rect -159 -1026 -129 -1000
rect -63 -1022 -33 -1000
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -273 -1088 -207 -1072
rect -81 -1038 -15 -1022
rect 33 -1026 63 -1000
rect 129 -1022 159 -1000
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect -81 -1088 -15 -1072
rect 111 -1038 177 -1022
rect 225 -1026 255 -1000
rect 321 -1022 351 -1000
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect 111 -1088 177 -1072
rect 303 -1038 369 -1022
rect 417 -1026 447 -1000
rect 513 -1022 543 -1000
rect 303 -1072 319 -1038
rect 353 -1072 369 -1038
rect 303 -1088 369 -1072
rect 495 -1038 561 -1022
rect 609 -1026 639 -1000
rect 705 -1022 735 -1000
rect 495 -1072 511 -1038
rect 545 -1072 561 -1038
rect 495 -1088 561 -1072
rect 687 -1038 753 -1022
rect 801 -1026 831 -1000
rect 897 -1022 927 -1000
rect 687 -1072 703 -1038
rect 737 -1072 753 -1038
rect 687 -1088 753 -1072
rect 879 -1038 945 -1022
rect 993 -1026 1023 -1000
rect 879 -1072 895 -1038
rect 929 -1072 945 -1038
rect 879 -1088 945 -1072
<< polycont >>
rect -929 1038 -895 1072
rect -737 1038 -703 1072
rect -545 1038 -511 1072
rect -353 1038 -319 1072
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect 415 1038 449 1072
rect 607 1038 641 1072
rect 799 1038 833 1072
rect 991 1038 1025 1072
rect -1025 -1072 -991 -1038
rect -833 -1072 -799 -1038
rect -641 -1072 -607 -1038
rect -449 -1072 -415 -1038
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
rect 319 -1072 353 -1038
rect 511 -1072 545 -1038
rect 703 -1072 737 -1038
rect 895 -1072 929 -1038
<< locali >>
rect -1187 1140 -1091 1174
rect 1091 1140 1187 1174
rect -1187 1078 -1153 1140
rect 1153 1078 1187 1140
rect -945 1038 -929 1072
rect -895 1038 -879 1072
rect -753 1038 -737 1072
rect -703 1038 -687 1072
rect -561 1038 -545 1072
rect -511 1038 -495 1072
rect -369 1038 -353 1072
rect -319 1038 -303 1072
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect 15 1038 31 1072
rect 65 1038 81 1072
rect 207 1038 223 1072
rect 257 1038 273 1072
rect 399 1038 415 1072
rect 449 1038 465 1072
rect 591 1038 607 1072
rect 641 1038 657 1072
rect 783 1038 799 1072
rect 833 1038 849 1072
rect 975 1038 991 1072
rect 1025 1038 1041 1072
rect -1073 988 -1039 1004
rect -1073 -1004 -1039 -988
rect -977 988 -943 1004
rect -977 -1004 -943 -988
rect -881 988 -847 1004
rect -881 -1004 -847 -988
rect -785 988 -751 1004
rect -785 -1004 -751 -988
rect -689 988 -655 1004
rect -689 -1004 -655 -988
rect -593 988 -559 1004
rect -593 -1004 -559 -988
rect -497 988 -463 1004
rect -497 -1004 -463 -988
rect -401 988 -367 1004
rect -401 -1004 -367 -988
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect 367 988 401 1004
rect 367 -1004 401 -988
rect 463 988 497 1004
rect 463 -1004 497 -988
rect 559 988 593 1004
rect 559 -1004 593 -988
rect 655 988 689 1004
rect 655 -1004 689 -988
rect 751 988 785 1004
rect 751 -1004 785 -988
rect 847 988 881 1004
rect 847 -1004 881 -988
rect 943 988 977 1004
rect 943 -1004 977 -988
rect 1039 988 1073 1004
rect 1039 -1004 1073 -988
rect -1041 -1072 -1025 -1038
rect -991 -1072 -975 -1038
rect -849 -1072 -833 -1038
rect -799 -1072 -783 -1038
rect -657 -1072 -641 -1038
rect -607 -1072 -591 -1038
rect -465 -1072 -449 -1038
rect -415 -1072 -399 -1038
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect 303 -1072 319 -1038
rect 353 -1072 369 -1038
rect 495 -1072 511 -1038
rect 545 -1072 561 -1038
rect 687 -1072 703 -1038
rect 737 -1072 753 -1038
rect 879 -1072 895 -1038
rect 929 -1072 945 -1038
rect -1187 -1140 -1153 -1078
rect 1153 -1140 1187 -1078
rect -1187 -1174 -1091 -1140
rect 1091 -1174 1187 -1140
<< viali >>
rect -929 1038 -895 1072
rect -737 1038 -703 1072
rect -545 1038 -511 1072
rect -353 1038 -319 1072
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect 415 1038 449 1072
rect 607 1038 641 1072
rect 799 1038 833 1072
rect 991 1038 1025 1072
rect -1073 -988 -1039 988
rect -977 -988 -943 988
rect -881 -988 -847 988
rect -785 -988 -751 988
rect -689 -988 -655 988
rect -593 -988 -559 988
rect -497 -988 -463 988
rect -401 -988 -367 988
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect 367 -988 401 988
rect 463 -988 497 988
rect 559 -988 593 988
rect 655 -988 689 988
rect 751 -988 785 988
rect 847 -988 881 988
rect 943 -988 977 988
rect 1039 -988 1073 988
rect -1025 -1072 -991 -1038
rect -833 -1072 -799 -1038
rect -641 -1072 -607 -1038
rect -449 -1072 -415 -1038
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
rect 319 -1072 353 -1038
rect 511 -1072 545 -1038
rect 703 -1072 737 -1038
rect 895 -1072 929 -1038
<< metal1 >>
rect -941 1072 -883 1078
rect -941 1038 -929 1072
rect -895 1038 -883 1072
rect -941 1032 -883 1038
rect -749 1072 -691 1078
rect -749 1038 -737 1072
rect -703 1038 -691 1072
rect -749 1032 -691 1038
rect -557 1072 -499 1078
rect -557 1038 -545 1072
rect -511 1038 -499 1072
rect -557 1032 -499 1038
rect -365 1072 -307 1078
rect -365 1038 -353 1072
rect -319 1038 -307 1072
rect -365 1032 -307 1038
rect -173 1072 -115 1078
rect -173 1038 -161 1072
rect -127 1038 -115 1072
rect -173 1032 -115 1038
rect 19 1072 77 1078
rect 19 1038 31 1072
rect 65 1038 77 1072
rect 19 1032 77 1038
rect 211 1072 269 1078
rect 211 1038 223 1072
rect 257 1038 269 1072
rect 211 1032 269 1038
rect 403 1072 461 1078
rect 403 1038 415 1072
rect 449 1038 461 1072
rect 403 1032 461 1038
rect 595 1072 653 1078
rect 595 1038 607 1072
rect 641 1038 653 1072
rect 595 1032 653 1038
rect 787 1072 845 1078
rect 787 1038 799 1072
rect 833 1038 845 1072
rect 787 1032 845 1038
rect 979 1072 1037 1078
rect 979 1038 991 1072
rect 1025 1038 1037 1072
rect 979 1032 1037 1038
rect -1079 988 -1033 1000
rect -1079 -988 -1073 988
rect -1039 -988 -1033 988
rect -1079 -1000 -1033 -988
rect -983 988 -937 1000
rect -983 -988 -977 988
rect -943 -988 -937 988
rect -983 -1000 -937 -988
rect -887 988 -841 1000
rect -887 -988 -881 988
rect -847 -988 -841 988
rect -887 -1000 -841 -988
rect -791 988 -745 1000
rect -791 -988 -785 988
rect -751 -988 -745 988
rect -791 -1000 -745 -988
rect -695 988 -649 1000
rect -695 -988 -689 988
rect -655 -988 -649 988
rect -695 -1000 -649 -988
rect -599 988 -553 1000
rect -599 -988 -593 988
rect -559 -988 -553 988
rect -599 -1000 -553 -988
rect -503 988 -457 1000
rect -503 -988 -497 988
rect -463 -988 -457 988
rect -503 -1000 -457 -988
rect -407 988 -361 1000
rect -407 -988 -401 988
rect -367 -988 -361 988
rect -407 -1000 -361 -988
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect 361 988 407 1000
rect 361 -988 367 988
rect 401 -988 407 988
rect 361 -1000 407 -988
rect 457 988 503 1000
rect 457 -988 463 988
rect 497 -988 503 988
rect 457 -1000 503 -988
rect 553 988 599 1000
rect 553 -988 559 988
rect 593 -988 599 988
rect 553 -1000 599 -988
rect 649 988 695 1000
rect 649 -988 655 988
rect 689 -988 695 988
rect 649 -1000 695 -988
rect 745 988 791 1000
rect 745 -988 751 988
rect 785 -988 791 988
rect 745 -1000 791 -988
rect 841 988 887 1000
rect 841 -988 847 988
rect 881 -988 887 988
rect 841 -1000 887 -988
rect 937 988 983 1000
rect 937 -988 943 988
rect 977 -988 983 988
rect 937 -1000 983 -988
rect 1033 988 1079 1000
rect 1033 -988 1039 988
rect 1073 -988 1079 988
rect 1033 -1000 1079 -988
rect -1037 -1038 -979 -1032
rect -1037 -1072 -1025 -1038
rect -991 -1072 -979 -1038
rect -1037 -1078 -979 -1072
rect -845 -1038 -787 -1032
rect -845 -1072 -833 -1038
rect -799 -1072 -787 -1038
rect -845 -1078 -787 -1072
rect -653 -1038 -595 -1032
rect -653 -1072 -641 -1038
rect -607 -1072 -595 -1038
rect -653 -1078 -595 -1072
rect -461 -1038 -403 -1032
rect -461 -1072 -449 -1038
rect -415 -1072 -403 -1038
rect -461 -1078 -403 -1072
rect -269 -1038 -211 -1032
rect -269 -1072 -257 -1038
rect -223 -1072 -211 -1038
rect -269 -1078 -211 -1072
rect -77 -1038 -19 -1032
rect -77 -1072 -65 -1038
rect -31 -1072 -19 -1038
rect -77 -1078 -19 -1072
rect 115 -1038 173 -1032
rect 115 -1072 127 -1038
rect 161 -1072 173 -1038
rect 115 -1078 173 -1072
rect 307 -1038 365 -1032
rect 307 -1072 319 -1038
rect 353 -1072 365 -1038
rect 307 -1078 365 -1072
rect 499 -1038 557 -1032
rect 499 -1072 511 -1038
rect 545 -1072 557 -1038
rect 499 -1078 557 -1072
rect 691 -1038 749 -1032
rect 691 -1072 703 -1038
rect 737 -1072 749 -1038
rect 691 -1078 749 -1072
rect 883 -1038 941 -1032
rect 883 -1072 895 -1038
rect 929 -1072 941 -1038
rect 883 -1078 941 -1072
<< properties >>
string FIXED_BBOX -1170 -1157 1170 1157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 22 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
