* NGSPICE file created from interdigitezed_exmaple.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_V4M8MU a_n73_n1000# a_15_n1000# a_n15_n1026# VSUBS
X0 a_15_n1000# a_n15_n1026# a_n73_n1000# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=150000u
.ends


* Top level circuit interdigitezed_exmaple

Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_40 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_41 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_30 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_42 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_43 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_31 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_32 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_20 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_21 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_10 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_44 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_33 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_22 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_11 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_45 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_34 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_23 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_12 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_35 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_24 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_13 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_36 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_25 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_14 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_37 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_26 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_15 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_38 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_27 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_16 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_39 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_28 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_17 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_29 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_18 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_19 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_0 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_1 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_3 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_2 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_4 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_5 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_6 VSS Drain2 VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_7 Drain2 VSS VSI1 VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_8 VSS Drain1 VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
Xsky130_fd_pr__nfet_01v8_lvt_V4M8MU_9 Drain1 VSS VRF VSS sky130_fd_pr__nfet_01v8_lvt_V4M8MU
.end

